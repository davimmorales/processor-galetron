module BIOS(clock, address, output_bios);
	 input [9:0] address;
	 input clock;
	 output [31:0] output_bios;
	 integer firstClock = 0;
	 reg [31:0] bios[28:0];

	 
	 always @ ( posedge clock ) begin
	 	 if (firstClock==0) begin

bios[0] <= 32'b01101100000000000000000000000000;//Nop
bios[1] <= 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
bios[2] <= 32'b01101010110000000000000000000101;//Loadi #5, #0 to r[22]
bios[3] <= 32'b01101010111000000000000000000110;//Loadi #6, #0 to r[23]
bios[4] <= 32'b01101011000000000000000000000111;//Loadi #7, #0 to r[24]
bios[5] <= 32'b01101011001000000000000000001000;//Loadi #8, #0 to r[25]
bios[6] <= 32'b10010101000101100000000000000000;//LoadHD m[r[22]] to r[8]
bios[7] <= 32'b10010101001101110000000000000000;//LoadHD m[r[23]] to r[9]
bios[8] <= 32'b10010101010110000000000000000000;//LoadHD m[r[24]] to r[10]
bios[9] <= 32'b10010101011110010000000000000000;//LoadHD m[r[25]] to r[11]
bios[10] <= 32'b01101000010000000000000000001111;//Loadi #15 to r[2]
bios[11] <= 32'b01101000011000000000000001000100;//Loadi #68 to r[3]
bios[12] <= 32'b01101000101000000000000000010101;//Loadi #21 to r[5]
bios[13] <= 32'b10000001000000000000000000000000;//Output r[8]
bios[14] <= 32'b10000001001000000000000000000000;//Output r[9]
bios[15] <= 32'b10000001010000000000000000000000;//Output r[10]
bios[16] <= 32'b10000001011000000000000000000000;//Output r[11]
bios[17] <= 32'b01101010000000000000000000000000;//Loadi #0 to r[16]
bios[18] <= 32'b01101010001000000000000000000001;//Loadi #1 to r[17]
bios[19] <= 32'b01101010010000000000000000000010;//Loadi #2 to r[18]
bios[20] <= 32'b10011100000000000000000000000000;//Nop
   
	 	 firstClock <= 1;
	 	 end
	 end
	 
	 assign output_bios = bios[address];
endmodule // BIOS
