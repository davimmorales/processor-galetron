module BIOS(address, output_bios);
	 input [11:0] address;
	 output [31:0] output_bios;
	 reg [31:0] bios[36:0];

initial begin

bios[0] = 32'b01101100000000000000000000000000;//Nop
bios[1] = 32'b01101000001000000001111110101001;//Loadi #8105 to r[1]
bios[2] = 32'b10000000001000000000000000000000;//Output r[1]
bios[3] <= 32'b01101100000000000000000000000000;//Nop
bios[4] = 32'b01100100001000000000000000000100;//Store r[1] in m[#4]
bios[5] = 32'b01100000010000000000000000000100;//Load m[#4] to r[2]
bios[6] <= 32'b01101100000000000000000000000000;//Nop
bios[7] = 32'b01101000001000000000100000000000;//Loadi #1, #0 to r[1]
bios[8] = 32'b10010100001000010000000000000000;//LoadHD m[r[1]] to r[1]
bios[9] <= 32'b01101100000000000000000000000000;//Nop
bios[10] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
bios[11] = 32'b01101000001000000000000000000000;//Loadi #0, #0 to r[1]
bios[12] = 32'b01101000010000000000000100000000;//Loadi #256 to r[2]
bios[13] = 32'b10010100011000010000000000000000;//LoadHD m[r[1]] to r[3]
bios[14] = 32'b01011100100000000001100000000000;//SLT if r[0] < r[3], r[4] = 1 else r[4] = 0
bios[15] = 32'b01111100000001000000000000000000;//Pre Branch r[4]
bios[16] = 32'b01001100000000000000000000000100;//Branch on Zero #4
bios[17] = 32'b10011000011000100000000000000000;//rStore r[3] in m[r[2]] 
bios[18] = 32'b00000100001000010000000000000001;//ADDi r[1], #1 to r[1]
bios[19] = 32'b00000100010000100000000000000001;//ADDi r[2], #1 to r[2]
bios[20] = 32'b01010100000000000000000000001101;//Jump to #13
bios[21] = 32'b01101000001000000000000000000000;//Loadi #0 to r[1]
bios[22] = 32'b01101000010000000000000100000000;//Loadi #256 to r[2]
bios[23] = 32'b01011100011000010001000000000000;//SLT if r[1] < r[2], r[3] = 1 else r[3] = 0
bios[24] = 32'b01111100000000110000000000000000;//Pre Branch r[3]
bios[25] = 32'b01001100000000000000000000000011;//Branch on Zero #3
bios[26] = 32'b10001000000000010000000000000000;//rStore r[0] in m[r[1]] 
bios[27] = 32'b00000100001000010000000000000001;//ADDi r[1], #1 to r[1]
bios[28] = 32'b01010100000000000000000000010111;//Jump to #23
bios[29] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
bios[30] = 32'b01101000001000000000000000000000;//Loadi #0 to r[1]
bios[31] = 32'b01101000010000000000000000000000;//Loadi #0 to r[2]
bios[32] = 32'b01101000011000000000000000000000;//Loadi #0 to r[3]
bios[33] = 32'b01101000100000000000000000000000;//Loadi #0 to r[4]
bios[34] = 32'b10011100000000000000000000000000;//Start Systemm
//	 	 bios[0] <= 32'b01101100000000000000000000000000;//Nop
//	 	 bios[1] <= 32'b01101001111000000100000000000000;//Loadi #1, #0 to r[15]
//	 	 bios[2] <= 32'b01110101100000000000000000000000;//Input to r[12]
//	 	 bios[3] <= 32'b10010001100011110000000000000000;//hdStore r[12] in m[r[15]] 
//	 	 bios[4] <= 32'b10010101000011110000000000000000;//LoadHD m[r[15]] to r[8]
//	 	 bios[5] <= 32'b10000001000000000000000000000000;//Output r[8]
//	 	 bios[6] <= 32'b01110000000000000000000000000000;//Hlt
		 end

	 
	 assign output_bios = bios[address];
endmodule // BIOS
