module BIOS(clock, address, output_bios);
	 input [9:0] address;
	 input clock;
	 output [31:0] output_bios;
	 integer firstClock = 0;
	 reg [31:0] bios[100:0];

	 
	 always @ ( posedge clock ) begin
	 	 if (firstClock==0) begin
	 	 bios[0] <= 32'b01101100000000000000000000000000;//Nop
	 	 bios[1] <= 32'b01110110101000000000000000000000;//Input to r[21]
	 	 bios[2] <= 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
	 	 bios[3] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 bios[4] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 bios[5] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 bios[6] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 bios[7] <= 32'b01001100000000000000000000010011;//Branch on Zero #19
	 	 bios[8] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 bios[9] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 bios[10] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 bios[11] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 bios[12] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 bios[13] <= 32'b01001100000000000000000000010000;//Branch on Zero #16
	 	 bios[14] <= 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
	 	 bios[15] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 bios[16] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 bios[17] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 bios[18] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 bios[19] <= 32'b01001100000000000000000000010111;//Branch on Zero #23
	 	 bios[20] <= 32'b01101010110000000000000000000011;//Loadi #3 to r[22]
	 	 bios[21] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 bios[22] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 bios[23] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 bios[24] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 bios[25] <= 32'b01001100000000000000000000001010;//Branch on Zero #10
	 	 bios[26] <= 32'b01010100000000000000000000100111;//Jump to #39
	 	 bios[27] <= 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
	 	 bios[28] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 bios[29] <= 32'b01010100000000000000000000000001;//Jump to #1
	 	 bios[30] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 bios[31] <= 32'b01101010110000000000001001100000;//Loadi #608 to r[22]
	 	 bios[32] <= 32'b10000110111101100000000000000000;//Loadr m[r[22]] to r[23]
	 	 bios[33] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 bios[34] <= 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
	 	 bios[35] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 bios[36] <= 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
	 	 bios[37] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 bios[38] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 bios[39] <= 32'b01010100000000000000000000000001;//Jump to #1
	 	 bios[40] <= 32'b10000010111000000000000000000000;//Output r[23]
	 	 bios[41] <= 32'b00000110110101100000000000000010;//ADDi r[22], #2 to r[22]
	 	 bios[42] <= 32'b01010100000000000000000000100000;//Jump to #32
	 	 bios[43] <= 32'b01110110101000000000000000000000;//Input to r[21]
	 	 bios[44] <= 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
	 	 bios[45] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 bios[46] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 bios[47] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 bios[48] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 bios[49] <= 32'b01001100000000000000000000001101;//Branch on Zero #13
	 	 bios[50] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 bios[51] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 bios[52] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 bios[53] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 bios[54] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 bios[55] <= 32'b01001100000000000000000000001011;//Branch on Zero #11
	 	 bios[56] <= 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
	 	 bios[57] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 bios[58] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 bios[59] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 bios[60] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 bios[61] <= 32'b01001100000000000000000000000100;//Branch on Zero #4
	 	 bios[62] <= 32'b01010100000000000000000001000110;//Jump to #70
	 	 bios[63] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 bios[64] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 bios[65] <= 32'b01010100000000000000000000101011;//Jump to #43
	 	 bios[66] <= 32'b01010100000000000000000000000001;//Jump to #1
	 	 bios[67] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 bios[68] <= 32'b01101010110000000100000000000000;//Loadi #1, #0 to r[22]
	 	 bios[69] <= 32'b10010110111101100000000000000000;//LoadHD m[r[22]] to r[23]
	 	 bios[70] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 bios[71] <= 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
	 	 bios[72] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 bios[73] <= 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
	 	 bios[74] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 bios[75] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 bios[76] <= 32'b01010100000000000000000000101011;//Jump to #43
	 	 bios[77] <= 32'b01101010101000000000000000000001;//Loadi #1 to r[21]
	 	 bios[78] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 bios[79] <= 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
	 	 bios[80] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 bios[81] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 bios[82] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 bios[83] <= 32'b10000010111000000000000000000000;//Output r[23]
	 	 bios[84] <= 32'b00000110110101100000000000100000;//ADDi r[22], #32 to r[22]
	 	 bios[85] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 bios[86] <= 32'b01010100000000000000000001000101;//Jump to #69
	 	 bios[87] <= 32'b01101010110000000000000111000010;//Loadi #450 to r[22]
	 	 bios[88] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 bios[89] <= 32'b01010100000000000000000000101011;//Jump to #43
	 	 bios[90] <= 32'b01101010110000000000000000000011;//Loadi #3 to r[22]
	 	 bios[91] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 bios[92] <= 32'b01010100000000000000000000000001;//Jump to #1
	 	 bios[93] <= 32'b01101010110000000000000111000010;//Loadi #450 to r[22]
	 	 bios[94] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 bios[95] <= 32'b01010100000000000000000000000001;//Jump to #1
	 	 bios[96] <= 32'b01010100000000000000000000000000;//Jump to #0
	 	 firstClock <= 1;
	 	 end
	 end
	 
	 assign output_bios = bios[address];
endmodule // BIOS
