module harddrive(data_write, track, sector, clock, output_hard_drive, flag_write_hd);
  input  [31:0] data_write;
  input [6:0] track;
  input [13:0] sector;
  input flag_write_hd;
  input clock;
  output [31:0] output_hard_drive;
  integer firstClock = 0;

	// Declare the hard drive variable
	reg [31:0] HD[1:0][1:0];

	always @ (posedge clock) begin
	//load instructions
	   if (firstClock==0) begin
//HD[1][0] <= 32'b00000000000000000000000000001001;
//HD[1][1] <= 32'b00000000000000000000000000000001;
//HD[1][2] <= 32'b00000000000000000000000000000000;
//HD[1][3] <= 32'b00000000000000000000000000000001;
//HD[1][32] <= 32'b00000000000000000000000000011111;
//HD[1][33] <= 32'b00000000000000000000000000000000;
//HD[1][34] <= 32'b00000000000000000000000000000001;
//HD[1][35] <= 32'b00000000000000000000000000000001;
//HD[1][64] <= 32'b00000000000000000000000000000100;
//HD[1][65] <= 32'b00000000000000000000000000000010;
//HD[1][66] <= 32'b00000000000000000000000000000001;
//HD[1][67] <= 32'b00000000000000000000000000000001;
//HD[1][96] <= 32'b00000000000000000000000000011000;
//HD[1][97] <= 32'b00000000000000000000000000001010;
//HD[1][98] <= 32'b00000000000000000000000000000001;
//HD[1][99] <= 32'b00000000000000000000000000000001;
//HD[1][128] <= 32'b00000000000000000000000000000000;
	//	HD[2][0] <= 32'b01101100000000000000000000000000;//Nop
	//	HD[2][1] <= 32'b01110101100000000000000000000000;//Input to r[12]
	//	HD[2][2] <= 32'b00000101100011000000000000000110;//ADDi r[12], #10 to r[12]
	//	HD[2][3] <= 32'b10000001100000000000000000000000;//Output r[12]
	//	HD[2][4] <= 32'b01110000000000000000000000000000;//Hlt
	//	HD[2][5] <= 32'b00000000000000000000000000000000;
	//	HD[2][24] <= 32'b01110100101000000000000000000000;//Input to r[5]
	 //	HD[2][25] <= 32'b00000100110001010000000000001010;//ADDi r[5], #10 to r[6]
	 //	HD[2][26] <= 32'b01100100110000000000000000001000;//Store r[6] in m[#8]
	 //	HD[2][27] <= 32'b01100001100000000000000000001000;//Load m[#8] to r[12]
	 //	HD[2][28] <= 32'b10000001100000000000000000000000;//Output r[12]
	 //	HD[2][29] <= 32'b01010100000000000000000000000111;//Jump to #7
	 //	HD[2][30] <= 32'b10000000101000000000000000000000;//Output r[5]
	 //	HD[2][31] <= 32'b01101001011000000000000110100100;//Loadi #420 to r[11]
	 //	HD[2][32] <= 32'b10000001011000000000000000000000;//Output r[11]
	//	HD[2][33] <= 32'b00000000000000000000000000000000;


			firstClock <= 1;
		end
	// Write
		if (flag_write_hd) begin
			HD[track][sector] <= data_write;
		end
	end


	// Continuous assignment implies read returns NEW data.
	// This is the natural behavior of the TriMatrix memory
	// blocks in Single Port mode.
	assign output_hard_drive = HD[track][sector];

endmodule
