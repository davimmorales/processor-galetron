module harddrive(data_write, hd_address, clock, output_hard_drive, flag_write_hd);
  input  [31:0] data_write;
  input [20:0] hd_address;
  input flag_write_hd;
  input clock;
  output [31:0] output_hard_drive;

	// Declare the hard drive variable
	reg [31:0] HD[12000:0];
   reg [20:0] hd_local_address;


	//operating system
	initial begin
  HD[0] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[1] = 32'b01110110101000000000000000000000;//Input to r[21]
  HD[2] = 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
  HD[3] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[4] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[5] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[6] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[7] = 32'b01001100000000000000000000010011;//Branch on Zero #19
  HD[8] = 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
  HD[9] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[10] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[11] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[12] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[13] = 32'b01001100000000000000000000010000;//Branch on Zero #16
  HD[14] = 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
  HD[15] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[16] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[17] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[18] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[19] = 32'b01001100000000000000000000010111;//Branch on Zero #23
  HD[20] = 32'b01101100000000000000000000000000;//Nop
  HD[21] = 32'b01101100000000000000000000000000;//Nop
  HD[22] = 32'b01101100000000000000000000000000;//Nop
  HD[23] = 32'b01101100000000000000000000000000;//Nop
  HD[24] = 32'b01101100000000000000000000000000;//Nop
  HD[25] = 32'b01101100000000000000000000000000;//Nop
  HD[26] = 32'b01010100000000000000001101010111;//Jump to #855
  HD[27] = 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
  HD[28] = 32'b10000010110000000000000000000000;//Output r[22]
  HD[29] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[30] = 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
  HD[31] = 32'b01101010110000000000000011000000;//Loadi #192 to r[22]
  HD[32] = 32'b10000110111101100000000000000000;//Loadr m[r[22]] to r[23]
  HD[33] = 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
  HD[34] = 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
  HD[35] = 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
  HD[36] = 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
  HD[37] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[38] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[39] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[40] = 32'b10000010111000000000000000000000;//Output r[23]
  HD[41] = 32'b00000110110101100000000000000010;//ADDi r[22], #2 to r[22]
  HD[42] = 32'b01010100000000000000000100100000;//Jump to #288
  HD[43] = 32'b01110110101000000000000000000000;//Input to r[21]
  HD[44] = 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
  HD[45] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[46] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[47] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[48] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[49] = 32'b01001100000000000000000000001101;//Branch on Zero #13
  HD[50] = 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
  HD[51] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[52] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[53] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[54] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[55] = 32'b01001100000000000000000000001011;//Branch on Zero #11
  HD[56] = 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
  HD[57] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[58] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[59] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[60] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[61] = 32'b01001100000000000000000000000100;//Branch on Zero #4
  HD[62] = 32'b01010100000000000000000101010111;//Jump to #343
  HD[63] = 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
  HD[64] = 32'b10000010110000000000000000000000;//Output r[22]
  HD[65] = 32'b01010100000000000000000100101011;//Jump to #299
  HD[66] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[67] = 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
  HD[68] = 32'b01101010110000000000100000000000;//Loadi #1, #0 to r[22]
  HD[69] = 32'b10010110111101100000000000000000;//LoadHD m[r[22]] to r[23]
  HD[70] = 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
  HD[71] = 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
  HD[72] = 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
  HD[73] = 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
  HD[74] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[75] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[76] = 32'b01010100000000000000000100101011;//Jump to #299
  HD[77] = 32'b01101010101000000000000000000001;//Loadi #1 to r[21]
  HD[78] = 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
  HD[79] = 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
  HD[80] = 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
  HD[81] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[82] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[83] = 32'b10000010111000000000000000000000;//Output r[23]
  HD[84] = 32'b00000110110101100000000000100000;//ADDi r[22], #32 to r[22]
  HD[85] = 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
  HD[86] = 32'b01010100000000000000000101000101;//Jump to #325
  HD[87] = 32'b01101010110000000000000000000011;//Loadi #3 to r[22]
  HD[88] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[89] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[90] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[91] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[92] = 32'b01001100000000000000000000000000;//Branch on Zero #0
  HD[93] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[94] = 32'b01101010110000000000000011000000;//Loadi #192 to r[22]
  HD[95] = 32'b10000110111101100000000000000000;//Loadr m[r[22]] to r[23]
  HD[96] = 32'b01011111000000001011100000000000;//SLT if r[0] < r[23], r[24] = 1 else r[24] = 0
  HD[97] = 32'b01011111001101110000000000000000;//SLT if r[23] < r[0], r[25] = 1 else r[25] = 0
  HD[98] = 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
  HD[99] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[100] = 32'b01001100000000000000000000001001;//Branch on Zero #9
  HD[101] = 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
  HD[102] = 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
  HD[103] = 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
  HD[104] = 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
  HD[105] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[106] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[107] = 32'b01010100000000000000000100101011;//Jump to #299
  HD[108] = 32'b00000110110101100000000000000010;//ADDi r[22], #2 to r[22]
  HD[109] = 32'b01010100000000000000000101011111;//Jump to #351
  HD[110] = 32'b01101010110000000000100000000000;//Loadi #1, #0 to r[22]
  HD[111] = 32'b10010110111101100000000000000000;//LoadHD m[r[22]] to r[23]
  HD[112] = 32'b01011111000000001011100000000000;//SLT if r[0] < r[23], r[24] = 1 else r[24] = 0
  HD[113] = 32'b01011111001101110000000000000000;//SLT if r[23] < r[0], r[25] = 1 else r[25] = 0
  HD[114] = 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
  HD[115] = 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
  HD[116] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[117] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[118] = 32'b01010100000000000000000100101011;//Jump to #299
  HD[119] = 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
  HD[120] = 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
  HD[121] = 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
  HD[122] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[123] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[124] = 32'b00000110110101100000000000100000;//ADDi r[22], #32 to r[22]
  HD[125] = 32'b01010100000000000000000101101111;//Jump to #367
  HD[126] = 32'b01100110101000000000000011101010;//Store r[21] in m[#234]
  HD[127] = 32'b01110110101000000000000000000000;//Input to r[21]
  HD[128] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[129] = 32'b01011110111101010000000000000000;//SLT if r[21] < r[0], r[23] = 1 else r[23] = 0
  HD[130] = 32'b01011111000000001010100000000000;//SLT if r[0] < r[21], r[24] = 1 else r[24] = 0
  HD[131] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[132] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[133] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[134] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[135] = 32'b01100010110000000000000011101010;//Load m[#234] to r[22]
  HD[136] = 32'b10000010110000000000000000000000;//Output r[22]
  HD[137] = 32'b01010100000000000000000101111111;//Jump to #383
  HD[138] = 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
  HD[139] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[140] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[141] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[142] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[143] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[144] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[145] = 32'b01010100000000000000000100101011;//Jump to #299
  HD[146] = 32'b01010100000000000000001001011110;//Jump to #606
  HD[147] = 32'b01101011011000000000001001000110;//Loadi #582 to r[27]
  HD[148] = 32'b01010100000000000000000110010101;//Jump to #405
  HD[149] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[150] = 32'b01100100000000000000000011100000;//Store r[0] in m[#224]
  HD[151] = 32'b01100100000000000000000011100010;//Store r[0] in m[#226]
  HD[152] = 32'b01101010101000000000000011000000;//Loadi #192 to r[21]
  HD[153] = 32'b01100110101000000000000011100011;//Store r[21] in m[#227]
  HD[154] = 32'b01100010101000000000000011100011;//Load m[#227] to r[21]
  HD[155] = 32'b10000110110101010000000000000000;//Loadr m[r[21]] to r[22]
  HD[156] = 32'b01011110111101100000000000000000;//SLT if r[22] < r[0], r[23] = 1 else r[23] = 0
  HD[157] = 32'b01011111000000001011000000000000;//SLT if r[0] < r[22], r[24] = 1 else r[24] = 0
  HD[158] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[159] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[160] = 32'b01001100000000000000000000010100;//Branch on Zero #20
  HD[161] = 32'b01101011000000000000000000000001;//Loadi #1 to r[24]
  HD[162] = 32'b01011111000110001011000000000000;//SLT if r[24] < r[22], r[24] = 1 else r[24] = 0
  HD[163] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[164] = 32'b01001100000000000000000000001100;//Branch on Zero #12
  HD[165] = 32'b01100010101000000000000011100011;//Load m[#227] to r[21]
  HD[166] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[167] = 32'b10000110110101010000000000000000;//Loadr m[r[21]] to r[22]
  HD[168] = 32'b01011110111101100000000000000000;//SLT if r[22] < r[0], r[23] = 1 else r[23] = 0
  HD[169] = 32'b01011111000000001011000000000000;//SLT if r[0] < r[22], r[24] = 1 else r[24] = 0
  HD[170] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[171] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[172] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[173] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[174] = 32'b01100011000000000000000011100010;//Load m[#226] to r[24]
  HD[175] = 32'b00000111000110000000000000000001;//ADDi r[24], #1 to r[24]
  HD[176] = 32'b01100111000000000000000011100010;//Store r[24] in m[#226]
  HD[177] = 32'b01100010101000000000000011100011;//Load m[#227] to r[21]
  HD[178] = 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
  HD[179] = 32'b01100110101000000000000011100011;//Store r[21] in m[#227]
  HD[180] = 32'b01010100000000000000000110011010;//Jump to #410
  HD[181] = 32'b01100010101000000000000011100010;//Load m[#226] to r[21]
  HD[182] = 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
  HD[183] = 32'b01011110110101101010100000000000;//SLT if r[22] < r[21], r[22] = 1 else r[22] = 0
  HD[184] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[185] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[186] = 32'b01101010101000000000000000000001;//Loadi #1 to r[21]
  HD[187] = 32'b01100110101000000000000011100000;//Store r[21] in m[#224]
  HD[188] = 32'b01101100000000000000000000000000;//Nop
  HD[189] = 32'b01101100000000000000000000000000;//Nop
  HD[190] = 32'b01101100000000000000000000000000;//Nop
  HD[191] = 32'b01101100000000000000000000000000;//Nop
  HD[192] = 32'b01101100000000000000000000000000;//Nop
  HD[193] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[194] = 32'b01100010101000000000000011101010;//Load m[#234] to r[21]
  HD[195] = 32'b01100110101000000000000100001111;//Store r[21] in m[#271]
  HD[196] = 32'b01101011011000000000000111110000;//Loadi #496 to r[27]
  HD[197] = 32'b01100010101000000000000011101010;//Load m[#234] to r[21]
  HD[198] = 32'b01100110101000000000000011100100;//Store r[21] in m[#228]
  HD[199] = 32'b01100100000000000000000011100101;//Store r[0] in m[#229]
  HD[200] = 32'b01100100000000000000000011100110;//Store r[0] in m[#230]
  HD[201] = 32'b01101010101000000000000000000001;//Loadi #1 to r[21]
  HD[202] = 32'b01100110101000000000000011100111;//Store r[21] in m[#231]
  HD[203] = 32'b01100100000000000000000011101000;//Store r[0] in m[#232]
  HD[204] = 32'b01100011110000000000000100001111;//Load m[#271] to r[30]
  HD[205] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[206] = 32'b01100110101000000000000011101001;//Store r[21] in m[#233]
  HD[207] = 32'b01100010101000000000000011101001;//Load m[#233] to r[21]
  HD[208] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[209] = 32'b01100010111000000000000011100100;//Load m[#228] to r[23]
  HD[210] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[211] = 32'b01011111001101111011000000000000;//SLT if r[23] < r[22], r[25] = 1 else r[25] = 0
  HD[212] = 32'b00100111000110001100100000000000;//OR r[24],r[25] to r[24]
  HD[213] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[214] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[215] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[216] = 32'b01010100000000000000000111001110;//Jump to #462
  HD[217] = 32'b01100010101000000000000011101001;//Load m[#233] to r[21]
  HD[218] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[219] = 32'b01100010110000000000000011100101;//Load m[#229] to r[22]
  HD[220] = 32'b10010010110101010000000000000000;//hdStore r[22] in m[r[21]]
  HD[221] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[222] = 32'b01100010110000000000000011100110;//Load m[#230] to r[22]
  HD[223] = 32'b10010010110101010000000000000000;//hdStore r[22] in m[r[21]]
  HD[224] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[225] = 32'b01100010110000000000000011100111;//Load m[#231] to r[22]
  HD[226] = 32'b10010010110101010000000000000000;//hdStore r[22] in m[r[21]]
  HD[227] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[228] = 32'b01100010110000000000000011101000;//Load m[#232] to r[22]
  HD[229] = 32'b10010010110101010000000000000000;//hdStore r[22] in m[r[21]]
  HD[230] = 32'b01101100000000000000000000000000;//Nop
  HD[231] = 32'b01101100000000000000000000000000;//Nop
  HD[232] = 32'b01101100000000000000000000000000;//Nop
  HD[233] = 32'b01101100000000000000000000000000;//Nop
  HD[234] = 32'b01101100000000000000000000000000;//Nop
  HD[235] = 32'b01101100000000000000000000000000;//Nop
  HD[236] = 32'b01101100000000000000000000000000;//Nop
  HD[237] = 32'b01101100000000000000000000000000;//Nop
  HD[238] = 32'b01101100000000000000000000000000;//Nop
  HD[239] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[240] = 32'b01101011011000000000001000001110;//Loadi #526 to r[27]
  HD[241] = 32'b01100010101000000000000011101010;//Load m[#234] to r[21]
  HD[242] = 32'b01100110101000000000000011101011;//Store r[21] in m[#235]
  HD[243] = 32'b01100100000000000000000011101100;//Store r[0] in m[#236]
  HD[244] = 32'b01010100000000000000000111110101;//Jump to #501
  HD[245] = 32'b01101010101000000000000011000000;//Loadi #192 to r[21]
  HD[246] = 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
  HD[247] = 32'b10000111000101010000000000000000;//Loadr m[r[21]] to r[24]
  HD[248] = 32'b01011110111101101100000000000000;//SLT if r[22] < r[24], r[23] = 1 else r[23] = 0
  HD[249] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[250] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[251] = 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
  HD[252] = 32'b01010100000000000000000111110111;//Jump to #503
  HD[253] = 32'b01100010110000000000000011101011;//Load m[#235] to r[22]
  HD[254] = 32'b01100010111000000000000011101100;//Load m[#236] to r[23]
  HD[255] = 32'b10001010110101010000000000000000;//rStore r[22] in m[r[21]]
  HD[256] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[257] = 32'b10001010111101010000000000000000;//rStore r[23] in m[r[21]]
  HD[258] = 32'b01101100000000000000000000000000;//Nop
  HD[259] = 32'b01101100000000000000000000000000;//Nop
  HD[260] = 32'b01101100000000000000000000000000;//Nop
  HD[261] = 32'b01101100000000000000000000000000;//Nop
  HD[262] = 32'b01101100000000000000000000000000;//Nop
  HD[263] = 32'b01101100000000000000000000000000;//Nop
  HD[264] = 32'b01101100000000000000000000000000;//Nop
  HD[265] = 32'b01101100000000000000000000000000;//Nop
  HD[266] = 32'b01101100000000000000000000000000;//Nop
  HD[267] = 32'b01101100000000000000000000000000;//Nop
  HD[268] = 32'b01101100000000000000000000000000;//Nop
  HD[269] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[270] = 32'b01100010101000000000000011101010;//Load m[#234] to r[21]
  HD[271] = 32'b01100110101000000000000011110001;//Store r[21] in m[#241]
  HD[272] = 32'b01101011011000000000001000101011;//Loadi #555 to r[27]
  HD[273] = 32'b01101100000000000000000000000000;//Nop
  HD[274] = 32'b01101010110000000000100000000000;//Loadi #1, #0 to r[22]
  HD[275] = 32'b01100110110000000000000011110011;//Store r[22] in m[#243]
  HD[276] = 32'b01100010101000000000000011110011;//Load m[#243] to r[21]
  HD[277] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[278] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[279] = 32'b01011111000101100000000000000000;//SLT if r[22] < r[0], r[24] = 1 else r[24] = 0
  HD[280] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[281] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[282] = 32'b01001100000000000000000000001110;//Branch on Zero #14
  HD[283] = 32'b01100011001000000000000011110001;//Load m[#241] to r[25]
  HD[284] = 32'b01011110111101101100100000000000;//SLT if r[22] < r[25], r[23] = 1 else r[23] = 0
  HD[285] = 32'b01011111000110011011000000000000;//SLT if r[25] < r[22], r[24] = 1 else r[24] = 0
  HD[286] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[287] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[288] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[289] = 32'b01001100000000000000000000000100;//Branch on Zero #4
  HD[290] = 32'b00000110110101010000000000000101;//ADDi r[21], #5 to r[22]
  HD[291] = 32'b10010110110101100000000000000000;//LoadHD m[r[22]] to r[22]
  HD[292] = 32'b01100110110000000000000011110010;//Store r[22] in m[#242]
  HD[293] = 32'b01010100000000000000001000101010;//Jump to #554
  HD[294] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[295] = 32'b01100110101000000000000011110011;//Store r[21] in m[#243]
  HD[296] = 32'b01010100000000000000001000010100;//Jump to #532
  HD[297] = 32'b01100100000000000000000011110010;//Store r[0] in m[#242]
  HD[298] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[299] = 32'b01100010101000000000000011110010;//Load m[#242] to r[21]
  HD[300] = 32'b01100110101000000000000011101110;//Store r[21] in m[#238]
  HD[301] = 32'b01101011011000000000001001000101;//Loadi #581 to r[27]
  HD[302] = 32'b01100100000000000000000011101111;//Store r[0] in m[#239]
  HD[303] = 32'b01101010101000000000000011000000;//Loadi #192 to r[21]
  HD[304] = 32'b01100010110000000000000011101110;//Load m[#238] to r[22]
  HD[305] = 32'b00010010101101011011000000000000;//TIMES r[21],r[22] to r[21]
  HD[306] = 32'b01101100000000000000000000000000;//Nop
  HD[307] = 32'b01101010110000000001000000000000;//Loadi #2, #0 to r[22]
  HD[308] = 32'b00000010101101011011000000000000;//ADD r[21],r[22] to r[21]
  HD[309] = 32'b01100110101000000000000011110000;//Store r[21] in m[#240]
  HD[310] = 32'b01100010101000000000000011110000;//Load m[#240] to r[21]
  HD[311] = 32'b01100010110000000000000011101111;//Load m[#239] to r[22]
  HD[312] = 32'b00000010101101011011000000000000;//ADD r[21],r[22] to r[21]
  HD[313] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[314] = 32'b01011110111101100000000000000000;//SLT if r[22] < r[0], r[23] = 1 else r[23] = 0
  HD[315] = 32'b01011111000000001011000000000000;//SLT if r[0] < r[22], r[24] = 1 else r[24] = 0
  HD[316] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[317] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[318] = 32'b01001100000000000000000000000101;//Branch on Zero #5
  HD[319] = 32'b01100010111000000000000011101111;//Load m[#239] to r[23]
  HD[320] = 32'b10011010110101110000000000000000;//rStore r[22] in m[r[23]]
  HD[321] = 32'b00000110111101110000000000000001;//ADDi r[23], #1 to r[23]
  HD[322] = 32'b01100110111000000000000011101111;//Store r[23] in m[#239]
  HD[323] = 32'b01010100000000000000001000110110;//Jump to #566
  HD[324] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[325] = 32'b01010100000000000000000000000000;//Jump to #0
  HD[326] = 32'b01101011011000000000001001010110;//Loadi #598 to r[27]
  HD[327] = 32'b01010100000000000000001001001000;//Jump to #584
  HD[328] = 32'b01100100000000000000000011110100;//Store r[0] in m[#244]
  HD[329] = 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
  HD[330] = 32'b01101010101000000000000011000000;//Loadi #192 to r[21]
  HD[331] = 32'b10000110111101010000000000000000;//Loadr m[r[21]] to r[23]
  HD[332] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[333] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[334] = 32'b01001100000000000000000000000100;//Branch on Zero #4
  HD[335] = 32'b01101011001000000000000000000001;//Loadi #1 to r[25]
  HD[336] = 32'b01100111001000000000000011110100;//Store r[25] in m[#244]
  HD[337] = 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
  HD[338] = 32'b01010100000000000000001001001011;//Jump to #587
  HD[339] = 32'b01101100000000000000000000000000;//Nop
  HD[340] = 32'b01101100000000000000000000000000;//Nop
  HD[341] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[342] = 32'b01100010101000000000000011110100;//Load m[#244] to r[21]
  HD[343] = 32'b01011110110101010000000000000000;//SLT if r[21] < r[0], r[22] = 1 else r[22] = 0
  HD[344] = 32'b01011110111000001010100000000000;//SLT if r[0] < r[21], r[23] = 1 else r[23] = 0
  HD[345] = 32'b00100110110101101011100000000000;//OR r[22],r[23] to r[22]
  HD[346] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[347] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[348] = 32'b01001100000000000000000000011011;//Branch on Zero #27
  HD[349] = 32'b01010100000000000000000111000010;//Jump to #450
  HD[350] = 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
  HD[351] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[352] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[353] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[354] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[355] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[356] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[357] = 32'b01010100000000000000001001000110;//Jump to #582
  HD[358] = 32'b01101010110000000000000000000011;//Loadi #3 to r[22]
  HD[359] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[360] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[361] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[362] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[363] = 32'b01001100000000000000001011110010;//Branch on Zero #754
  HD[364] = 32'b01101010110000000000000000000100;//Loadi #4 to r[22]
  HD[365] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[366] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[367] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[368] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[369] = 32'b01001100000000000000000000000000;//Branch on Zero #0
  HD[370] = 32'b01101010110000000000000000000101;//Loadi #5 to r[22]
  HD[371] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[372] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[373] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[374] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[375] = 32'b01001100000000000000000000000000;//Branch on Zero #0
  HD[376] = 32'b01101011011000000000001001111010;//Loadi #634 to r[27]
  HD[377] = 32'b01101100000000000000000000000000;//Nop
  HD[378] = 32'b01101100000000000000000000000000;//Nop
  HD[379] = 32'b01101100000000000000000000000000;//Nop
  HD[380] = 32'b01101100000000000000000000000000;//Nop
  HD[381] = 32'b01101100000000000000000000000000;//Nop
  HD[382] = 32'b01101100000000000000000000000000;//Nop
  HD[383] = 32'b01101100000000000000000000000000;//Nop
  HD[384] = 32'b01101100000000000000000000000000;//Nop
  HD[385] = 32'b01101100000000000000000000000000;//Nop
  HD[386] = 32'b01101011011000000000001010100110;//Loadi #678 to r[27]
  HD[387] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[388] = 32'b01100110101000000000000011110110;//Store r[21] in m[#246]
  HD[389] = 32'b01100010101000000000000011110110;//Load m[#246] to r[21]
  HD[390] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[391] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[392] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[393] = 32'b01001100000000000000000000010100;//Branch on Zero #20
  HD[394] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[395] = 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
  HD[396] = 32'b01011111001000001011100000000000;//SLT if r[0] < r[23], r[25] = 1 else r[25] = 0
  HD[397] = 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
  HD[398] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[399] = 32'b01001100000000000000000000001011;//Branch on Zero #11
  HD[400] = 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
  HD[401] = 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
  HD[402] = 32'b01101011000000000000000000000001;//Loadi #1 to r[24]
  HD[403] = 32'b01011111001110001011100000000000;//SLT if r[24] < r[23], r[25] = 1 else r[25] = 0
  HD[404] = 32'b01011111000101111100000000000000;//SLT if r[23] < r[24], r[24] = 1 else r[24] = 0
  HD[405] = 32'b00100111001110011100000000000000;//OR r[25],r[24] to r[25]
  HD[406] = 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
  HD[407] = 32'b01111100000110010000000000000000;//Pre Branch r[25]
  HD[408] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[409] = 32'b01100110110000000000000011110111;//Store r[22] in m[#247]
  HD[410] = 32'b01010100000000000000001010011110;//Jump to #670
  HD[411] = 32'b01100010101000000000000011110110;//Load m[#246] to r[21]
  HD[412] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[413] = 32'b01010100000000000000001010000100;//Jump to #644
  HD[414] = 32'b01101100000000000000000000000000;//Nop
  HD[415] = 32'b01101100000000000000000000000000;//Nop
  HD[416] = 32'b01101100000000000000000000000000;//Nop
  HD[417] = 32'b01101100000000000000000000000000;//Nop
  HD[418] = 32'b01101100000000000000000000000000;//Nop
  HD[419] = 32'b01101100000000000000000000000000;//Nop
  HD[420] = 32'b01101100000000000000000000000000;//Nop
  HD[421] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[422] = 32'b01101011011000000000001011100001;//Loadi #737 to r[27]
  HD[423] = 32'b01101100000000000000000000000000;//Nop
  HD[424] = 32'b01101010101000000000000000000011;//Loadi #3 to r[21]
  HD[425] = 32'b01100110101000000000000011111001;//Store r[21] in m[#249]
  HD[426] = 32'b01100100000000000000000100001010;//Store r[0] in m[#266]
  HD[427] = 32'b01100100000000000000000100001011;//Store r[0] in m[#267]
  HD[428] = 32'b01100100000000000000000100001100;//Store r[0] in m[#268]
  HD[429] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[430] = 32'b01100110101000000000000011111000;//Store r[21] in m[#248]
  HD[431] = 32'b01100010101000000000000011111000;//Load m[#248] to r[21]
  HD[432] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[433] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[434] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[435] = 32'b01001100000000000000000000010100;//Branch on Zero #20
  HD[436] = 32'b01101010111000000000000000000001;//Loadi #1 to r[23]
  HD[437] = 32'b01011111000101111011000000000000;//SLT if r[23] < r[22], r[24] = 1 else r[24] = 0
  HD[438] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[439] = 32'b01001100000000000000000000001101;//Branch on Zero #13
  HD[440] = 32'b00000110101101010000000000000011;//ADDi r[21], #3 to r[21]
  HD[441] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[442] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[443] = 32'b01101100000000000000000000000000;//Nop
  HD[444] = 32'b01101100000000000000000000000000;//Nop
  HD[445] = 32'b00110111000110000000000000000000;//NOT r[24] to r[24]
  HD[446] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[447] = 32'b01001100000000000000000000000101;//Branch on Zero #5
  HD[448] = 32'b00001110101101010000000000000010;//SUBi r[21], #2 to r[21]
  HD[449] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[450] = 32'b01101011000000000000000100001010;//Loadi #266 to r[24]
  HD[451] = 32'b00000010110101101100000000000000;//ADD r[22],r[24] to r[22]
  HD[452] = 32'b10001010111101100000000000000000;//rStore r[23] in m[r[22]]
  HD[453] = 32'b01100010101000000000000011111000;//Load m[#248] to r[21]
  HD[454] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[455] = 32'b01010100000000000000001010101110;//Jump to #686
  HD[456] = 32'b01100010101000000000000100001011;//Load m[#267] to r[21]
  HD[457] = 32'b01011110110000001010100000000000;//SLT if r[0] < r[21], r[22] = 1 else r[22] = 0
  HD[458] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[459] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[460] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[461] = 32'b01101010111000000000000000000001;//Loadi #1 to r[23]
  HD[462] = 32'b01100110111000000000000011111001;//Store r[23] in m[#249]
  HD[463] = 32'b01010100000000000000001011010111;//Jump to #727
  HD[464] = 32'b01100010101000000000000100001100;//Load m[#268] to r[21]
  HD[465] = 32'b01011110110000001010100000000000;//SLT if r[0] < r[21], r[22] = 1 else r[22] = 0
  HD[466] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[467] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[468] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[469] = 32'b01101010111000000000000000000010;//Loadi #2 to r[23]
  HD[470] = 32'b01100110111000000000000011111001;//Store r[23] in m[#249]
  HD[471] = 32'b01101100000000000000000000000000;//Nop
  HD[472] = 32'b01101100000000000000000000000000;//Nop
  HD[473] = 32'b01101100000000000000000000000000;//Nop
  HD[474] = 32'b01101100000000000000000000000000;//Nop
  HD[475] = 32'b01101100000000000000000000000000;//Nop
  HD[476] = 32'b01101100000000000000000000000000;//Nop
  HD[477] = 32'b01101100000000000000000000000000;//Nop
  HD[478] = 32'b01101100000000000000000000000000;//Nop
  HD[479] = 32'b01101100000000000000000000000000;//Nop
  HD[480] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[481] = 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
  HD[482] = 32'b01100110101000000000000011111010;//Store r[21] in m[#250]
  HD[483] = 32'b01100010101000000000000011111001;//Load m[#249] to r[21]
  HD[484] = 32'b01100110101000000000000011111011;//Store r[21] in m[#251]
  HD[485] = 32'b01101011011000000000001100010100;//Loadi #788 to r[27]
  HD[486] = 32'b01101100000000000000000000000000;//Nop
  HD[487] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[488] = 32'b01100110101000000000000011111100;//Store r[21] in m[#252]
  HD[489] = 32'b01100010101000000000000011111100;//Load m[#252] to r[21]
  HD[490] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[491] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[492] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[493] = 32'b01001100000000000000000000010000;//Branch on Zero #16
  HD[494] = 32'b01100010111000000000000011111010;//Load m[#250] to r[23]
  HD[495] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[496] = 32'b01011110111101111011000000000000;//SLT if r[23] < r[22], r[23] = 1 else r[23] = 0
  HD[497] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[498] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[499] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[500] = 32'b01001100000000000000000000000110;//Branch on Zero #6
  HD[501] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[502] = 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
  HD[503] = 32'b01100110111000000000000011111101;//Store r[23] in m[#253]
  HD[504] = 32'b01100010111000000000000011111011;//Load m[#251] to r[23]
  HD[505] = 32'b10010010111101010000000000000000;//hdStore r[23] in m[r[21]]
  HD[506] = 32'b01010100000000000000001011111110;//Jump to #766
  HD[507] = 32'b01100010101000000000000011111100;//Load m[#252] to r[21]
  HD[508] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[509] = 32'b01010100000000000000001011101000;//Jump to #744
  HD[510] = 32'b01100010110000000000000011111101;//Load m[#253] to r[22]
  HD[511] = 32'b01101010111000000000000000100110;//Loadi #38 to r[23]
  HD[512] = 32'b00010010110101101011100000000000;//TIMES r[22],r[23] to r[22]
  HD[513] = 32'b01100110110000000000000011111101;//Store r[22] in m[#253]
  HD[514] = 32'b01100010110000000000000011111011;//Load m[#251] to r[22]
  HD[515] = 32'b00010010110101101011100000000000;//TIMES r[22],r[23] to r[22]
  HD[516] = 32'b01100110110000000000000011111110;//Store r[22] in m[#254]
  HD[517] = 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
  HD[518] = 32'b01100110101000000000000011111100;//Store r[21] in m[#252]
  HD[519] = 32'b01100010101000000000000011111100;//Load m[#252] to r[21]
  HD[520] = 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
  HD[521] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[522] = 32'b01001100000000000000000000001000;//Branch on Zero #8
  HD[523] = 32'b01100010110000000000000011111101;//Load m[#253] to r[22]
  HD[524] = 32'b00000010110101011011000000000000;//ADD r[21],r[22] to r[22]
  HD[525] = 32'b10000110110101100000000000000000;//Loadr m[r[22]] to r[22]
  HD[526] = 32'b01100011000000000000000011111110;//Load m[#254] to r[24]
  HD[527] = 32'b00000011000101011100000000000000;//ADD r[21],r[24] to r[24]
  HD[528] = 32'b10001010110110000000000000000000;//rStore r[22] in m[r[24]]
  HD[529] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[530] = 32'b01010100000000000000001100000110;//Jump to #774
  HD[531] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[532] = 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
  HD[533] = 32'b01100110101000000000000011111111;//Store r[21] in m[#255]
  HD[534] = 32'b01101011011000000000000111000010;//Loadi #450 to r[27]
  HD[535] = 32'b10000010100000000000000000000000;//Output r[20]
  HD[536] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[537] = 32'b01100110101000000000000100000000;//Store r[21] in m[#256]
  HD[538] = 32'b01100010101000000000000100000000;//Load m[#256] to r[21]
  HD[539] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[540] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[541] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[542] = 32'b01001100000000000000000000001011;//Branch on Zero #11
  HD[543] = 32'b01100010111000000000000011111111;//Load m[#255] to r[23]
  HD[544] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[545] = 32'b01011111001101111011000000000000;//SLT if r[23] < r[22], r[25] = 1 else r[25] = 0
  HD[546] = 32'b00100111000110001100100000000000;//OR r[24],r[25] to r[24]
  HD[547] = 32'b00110111000110000000000000000000;//NOT r[24] to r[24]
  HD[548] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[549] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[550] = 32'b01010100000000000000001100101010;//Jump to #810
  HD[551] = 32'b01100010101000000000000100000000;//Load m[#256] to r[21]
  HD[552] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[553] = 32'b01010100000000000000001100011001;//Jump to #793
  HD[554] = 32'b01100110101000000000000100000000;//Store r[21] in m[#256]
  HD[555] = 32'b01100010101000000000000100000000;//Load m[#256] to r[21]
  HD[556] = 32'b00000110101101010000000000000100;//ADDi r[21], #4 to r[21]
  HD[557] = 32'b10010011100101010000000000000000;//hdStore r[28] in m[r[21]]
  HD[558] = 32'b00000110101101010000000000001000;//ADDi r[21], #8 to r[21]
  HD[559] = 32'b10010000000101010000000000000000;//hdStore r[0] in m[r[21]]
  HD[560] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[561] = 32'b10010000001101010000000000000000;//hdStore r[1] in m[r[21]]
  HD[562] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[563] = 32'b10010000010101010000000000000000;//hdStore r[2] in m[r[21]]
  HD[564] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[565] = 32'b10010000011101010000000000000000;//hdStore r[3] in m[r[21]]
  HD[566] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[567] = 32'b10010000100101010000000000000000;//hdStore r[4] in m[r[21]]
  HD[568] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[569] = 32'b10010000101101010000000000000000;//hdStore r[5] in m[r[21]]
  HD[570] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[571] = 32'b10010000110101010000000000000000;//hdStore r[6] in m[r[21]]
  HD[572] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[573] = 32'b10010000111101010000000000000000;//hdStore r[7] in m[r[21]]
  HD[574] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[575] = 32'b10010001000101010000000000000000;//hdStore r[8] in m[r[21]]
  HD[576] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[577] = 32'b10010001001101010000000000000000;//hdStore r[9] in m[r[21]]
  HD[578] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[579] = 32'b10010001010101010000000000000000;//hdStore r[10] in m[r[21]]
  HD[580] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[581] = 32'b10010001011101010000000000000000;//hdStore r[11] in m[r[21]]
  HD[582] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[583] = 32'b10010001100101010000000000000000;//hdStore r[12] in m[r[21]]
  HD[584] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[585] = 32'b10010001101101010000000000000000;//hdStore r[13] in m[r[21]]
  HD[586] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[587] = 32'b10010001110101010000000000000000;//hdStore r[14] in m[r[21]]
  HD[588] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[589] = 32'b10010001111101010000000000000000;//hdStore r[15] in m[r[21]]
  HD[590] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[591] = 32'b10010010000101010000000000000000;//hdStore r[16] in m[r[21]]
  HD[592] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[593] = 32'b10010010001101010000000000000000;//hdStore r[17] in m[r[21]]
  HD[594] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[595] = 32'b10010010010101010000000000000000;//hdStore r[18] in m[r[21]]
  HD[596] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[597] = 32'b10010010011101010000000000000000;//hdStore r[19] in m[r[21]]
  HD[598] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[599] = 32'b01101010110000000000000000001010;//Loadi #10 to r[22]
  HD[600] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[601] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[602] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[603] = 32'b01010100000000000000010011011101;//Jump to #1245
  HD[604] = 32'b01100110101000000000000100000100;//Store r[21] in m[#260]
  HD[605] = 32'b01100110101000000000000100000001;//Store r[21] in m[#257]
  HD[606] = 32'b01101011011000000000001101111111;//Loadi #895 to r[27]
  HD[607] = 32'b01010100000000000000001101100000;//Jump to #864
  HD[608] = 32'b01100100000000000000000100000011;//Store r[0] in m[#259]
  HD[609] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[610] = 32'b01100110101000000000000100000010;//Store r[21] in m[#258]
  HD[611] = 32'b01100010101000000000000100000010;//Load m[#258] to r[21]
  HD[612] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[613] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[614] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[615] = 32'b01001100000000000000000000010101;//Branch on Zero #21
  HD[616] = 32'b01100010111000000000000100000001;//Load m[#257] to r[23]
  HD[617] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[618] = 32'b01011110111101111011000000000000;//SLT if r[23] < r[22], r[23] = 1 else r[23] = 0
  HD[619] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[620] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[621] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[622] = 32'b01001100000000000000000000001011;//Branch on Zero #11
  HD[623] = 32'b00000110101101010000000000000011;//ADDi r[21], #3 to r[21]
  HD[624] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[625] = 32'b01101010111000000000000000000001;//Loadi #1 to r[23]
  HD[626] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[627] = 32'b01101100000000000000000000000000;//Nop
  HD[628] = 32'b01101100000000000000000000000000;//Nop
  HD[629] = 32'b00110111000110000000000000000000;//NOT r[24] to r[24]
  HD[630] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[631] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[632] = 32'b01100110111000000000000100000011;//Store r[23] in m[#259]
  HD[633] = 32'b01010100000000000000001101111101;//Jump to #893
  HD[634] = 32'b01100010101000000000000100000010;//Load m[#258] to r[21]
  HD[635] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[636] = 32'b01010100000000000000001101100010;//Jump to #866
  HD[637] = 32'b01101100000000000000000000000000;//Nop
  HD[638] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[639] = 32'b01100010101000000000000100000011;//Load m[#259] to r[21]
  HD[640] = 32'b01011110110000001010100000000000;//SLT if r[0] < r[21], r[22] = 1 else r[22] = 0
  HD[641] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[642] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[643] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[644] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[645] = 32'b01110110101000000000000000000000;//Input to r[21]
  HD[646] = 32'b01011110110000001010100000000000;//SLT if r[0] < r[21], r[22] = 1 else r[22] = 0
  HD[647] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[648] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[649] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[650] = 32'b01100010110000000000000100000100;//Load m[#260] to r[22]
  HD[651] = 32'b10000010110000000000000000000000;//Output r[22]
  HD[652] = 32'b01010100000000000000001110000101;//Jump to #901
  HD[653] = 32'b01101011000000000000000000000010;//Loadi #2 to r[24]
  HD[654] = 32'b01011110110101011100000000000000;//SLT if r[21] < r[24], r[22] = 1 else r[22] = 0
  HD[655] = 32'b01011110111110001010100000000000;//SLT if r[24] < r[21], r[23] = 1 else r[23] = 0
  HD[656] = 32'b00100110110101101011100000000000;//OR r[22],r[23] to r[22]
  HD[657] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[658] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[659] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[660] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[661] = 32'b01101011000000000000000000000011;//Loadi #3 to r[24]
  HD[662] = 32'b01011110110101011100000000000000;//SLT if r[21] < r[24], r[22] = 1 else r[22] = 0
  HD[663] = 32'b01011110111110001010100000000000;//SLT if r[24] < r[21], r[23] = 1 else r[23] = 0
  HD[664] = 32'b00100110110101101011100000000000;//OR r[22],r[23] to r[22]
  HD[665] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[666] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[667] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[668] = 32'b01010100000000000000010101001011;//Jump to #1355
  HD[669] = 32'b01011110110110001010100000000000;//SLT if r[24] < r[21], r[22] = 1 else r[22] = 0
  HD[670] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[671] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[672] = 32'b01010100000000000000001110000101;//Jump to #901
  HD[673] = 32'b01101011000000000000000000000001;//Loadi #1 to r[24]
  HD[674] = 32'b01011110110101011100000000000000;//SLT if r[21] < r[24], r[22] = 1 else r[22] = 0
  HD[675] = 32'b01011110111110001010100000000000;//SLT if r[24] < r[21], r[23] = 1 else r[23] = 0
  HD[676] = 32'b00100110110101101011100000000000;//OR r[22],r[23] to r[22]
  HD[677] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[678] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[679] = 32'b01010100000000000000001110000101;//Jump to #901
  HD[680] = 32'b01100010101000000000000100000100;//Load m[#260] to r[21]
  HD[681] = 32'b01100110101000000000000100000101;//Store r[21] in m[#261]
  HD[682] = 32'b01100110101000000000000100001111;//Store r[21] in m[#271]
  HD[683] = 32'b01101011011000000000010101000011;//Loadi #1347 to r[27]
  HD[684] = 32'b01100011110000000000000100001111;//Load m[#271] to r[30]
  HD[685] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[686] = 32'b01100110101000000000000100000110;//Store r[21] in m[#262]
  HD[687] = 32'b01100010101000000000000100000110;//Load m[#262] to r[21]
  HD[688] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[689] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[690] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[691] = 32'b01001100000000000000000000010100;//Branch on Zero #20
  HD[692] = 32'b01101011000000000000000000000001;//Loadi #1 to r[24]
  HD[693] = 32'b01011110111101101100000000000000;//SLT if r[22] < r[24], r[23] = 1 else r[23] = 0
  HD[694] = 32'b01011111000110001011000000000000;//SLT if r[24] < r[22], r[24] = 1 else r[24] = 0
  HD[695] = 32'b00100111000110001011100000000000;//OR r[24],r[23] to r[24]
  HD[696] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[697] = 32'b01001100000000000000000000001011;//Branch on Zero #11
  HD[698] = 32'b01100011000000000000000100000101;//Load m[#261] to r[24]
  HD[699] = 32'b01011110111101101100000000000000;//SLT if r[22] < r[24], r[23] = 1 else r[23] = 0
  HD[700] = 32'b01011111000110001011000000000000;//SLT if r[24] < r[22], r[24] = 1 else r[24] = 0
  HD[701] = 32'b00100111000110001011100000000000;//OR r[24],r[23] to r[24]
  HD[702] = 32'b00110111000110000000000000000000;//NOT r[24] to r[24]
  HD[703] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[704] = 32'b01001100000000000000000000000100;//Branch on Zero #4
  HD[705] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[706] = 32'b10010111000101010000000000000000;//LoadHD m[r[21]] to r[24]
  HD[707] = 32'b01100111000000000000000100000111;//Store r[24] in m[#263]
  HD[708] = 32'b01010100000000000000001111001000;//Jump to #968
  HD[709] = 32'b01100010101000000000000100000110;//Load m[#262] to r[21]
  HD[710] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[711] = 32'b01010100000000000000001110101110;//Jump to #942
  HD[712] = 32'b01101100000000000000000000000000;//Nop
  HD[713] = 32'b01101100000000000000000000000000;//Nop
  HD[714] = 32'b01101100000000000000000000000000;//Nop
  HD[715] = 32'b01101100000000000000000000000000;//Nop
  HD[716] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[717] = 32'b01100010101000000000000100000100;//Load m[#260] to r[21]
  HD[718] = 32'b01100110101000000000000011111010;//Store r[21] in m[#250]
  HD[719] = 32'b01101010101000000000000000000100;//Loadi #4 to r[21]
  HD[720] = 32'b01100110101000000000000011111011;//Store r[21] in m[#251]
  HD[721] = 32'b01101011011000000000001111010011;//Loadi #979 to r[27]
  HD[722] = 32'b01010100000000000000001011100111;//Jump to #743
  HD[723] = 32'b01101011011000000000001111010101;//Loadi #981 to r[27]
  HD[724] = 32'b01010100000000000000001010000011;//Jump to #643
  HD[725] = 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
  HD[726] = 32'b01100110101000000000000011111010;//Store r[21] in m[#250]
  HD[727] = 32'b01100010101000000000000100000111;//Load m[#263] to r[21]
  HD[728] = 32'b01100110101000000000000011111011;//Store r[21] in m[#251]
  HD[729] = 32'b01101011011000000000001111011011;//Loadi #987 to r[27]
  HD[730] = 32'b01010100000000000000001011100111;//Jump to #743
  HD[731] = 32'b01100010101000000000000100000100;//Load m[#260] to r[21]
  HD[732] = 32'b01100110101000000000000011111010;//Store r[21] in m[#250]
  HD[733] = 32'b01100100000000000000000011111011;//Store r[0] in m[#251]
  HD[734] = 32'b01101011011000000000001111100000;//Loadi #992 to r[27]
  HD[735] = 32'b01010100000000000000001011100111;//Jump to #743
  HD[736] = 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
  HD[737] = 32'b01100110101000000000000011111111;//Store r[21] in m[#255]
  HD[738] = 32'b01101011011000000000001111100100;//Loadi #996 to r[27]
  HD[739] = 32'b01010100000000000000001100011000;//Jump to #792
  HD[740] = 32'b01100010101000000000000100000100;//Load m[#260] to r[21]
  HD[741] = 32'b01100110101000000000000100001000;//Store r[21] in m[#264]
  HD[742] = 32'b01101011011000000000010000101011;//Loadi #1067 to r[27]
  HD[743] = 32'b01010100000000000000001111101000;//Jump to #1000
  HD[744] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[745] = 32'b01100110101000000000000100001001;//Store r[21] in m[#265]
  HD[746] = 32'b01100010101000000000000100001001;//Load m[#265] to r[21]
  HD[747] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[748] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[749] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[750] = 32'b01001100000000000000000000001011;//Branch on Zero #11
  HD[751] = 32'b01100010111000000000000100001000;//Load m[#264] to r[23]
  HD[752] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[753] = 32'b01011111001101111011000000000000;//SLT if r[23] < r[22], r[25] = 1 else r[25] = 0
  HD[754] = 32'b00100111000110001100100000000000;//OR r[24],r[25] to r[24]
  HD[755] = 32'b00110111000110000000000000000000;//NOT r[24] to r[24]
  HD[756] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[757] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[758] = 32'b01010100000000000000001111111010;//Jump to #1018
  HD[759] = 32'b01100010101000000000000100001001;//Load m[#265] to r[21]
  HD[760] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[761] = 32'b01010100000000000000001111101001;//Jump to #1001
  HD[762] = 32'b01100110101000000000000100001001;//Store r[21] in m[#265]
  HD[763] = 32'b01100010101000000000000100001001;//Load m[#265] to r[21]
  HD[764] = 32'b00000110101101010000000000000100;//ADDi r[21], #4 to r[21]
  HD[765] = 32'b10010111100101010000000000000000;//LoadHD m[r[21]] to r[28]
  HD[766] = 32'b00000110101101010000000000001000;//ADDi r[21], #8 to r[21]
  HD[767] = 32'b10010100000101010000000000000000;//LoadHD m[r[21]] to r[0]
  HD[768] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[769] = 32'b10010100001101010000000000000000;//LoadHD m[r[21]] to r[1]
  HD[770] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[771] = 32'b10010100010101010000000000000000;//LoadHD m[r[21]] to r[2]
  HD[772] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[773] = 32'b10010100011101010000000000000000;//LoadHD m[r[21]] to r[3]
  HD[774] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[775] = 32'b10010100100101010000000000000000;//LoadHD m[r[21]] to r[4]
  HD[776] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[777] = 32'b10010100101101010000000000000000;//LoadHD m[r[21]] to r[5]
  HD[778] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[779] = 32'b10010100110101010000000000000000;//LoadHD m[r[21]] to r[6]
  HD[780] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[781] = 32'b10010100111101010000000000000000;//LoadHD m[r[21]] to r[7]
  HD[782] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[783] = 32'b10010101000101010000000000000000;//LoadHD m[r[21]] to r[8]
  HD[784] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[785] = 32'b10010101001101010000000000000000;//LoadHD m[r[21]] to r[9]
  HD[786] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[787] = 32'b10010101010101010000000000000000;//LoadHD m[r[21]] to r[10]
  HD[788] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[789] = 32'b10010101011101010000000000000000;//LoadHD m[r[21]] to r[11]
  HD[790] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[791] = 32'b10010101100101010000000000000000;//LoadHD m[r[21]] to r[12]
  HD[792] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[793] = 32'b10010101101101010000000000000000;//LoadHD m[r[21]] to r[13]
  HD[794] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[795] = 32'b10010101110101010000000000000000;//LoadHD m[r[21]] to r[14]
  HD[796] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[797] = 32'b10010101111101010000000000000000;//LoadHD m[r[21]] to r[15]
  HD[798] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[799] = 32'b10010110000101010000000000000000;//LoadHD m[r[21]] to r[16]
  HD[800] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[801] = 32'b10010110001101010000000000000000;//LoadHD m[r[21]] to r[17]
  HD[802] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[803] = 32'b10010110010101010000000000000000;//LoadHD m[r[21]] to r[18]
  HD[804] = 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
  HD[805] = 32'b10010110011101010000000000000000;//LoadHD m[r[21]] to r[19]
  HD[806] = 32'b01101100000000000000000000000000;//Nop
  HD[807] = 32'b01101100000000000000000000000000;//Nop
  HD[808] = 32'b01101100000000000000000000000000;//Nop
  HD[809] = 32'b01101100000000000000000000000000;//Nop
  HD[810] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[811] = 32'b01101011011000000000010000101111;//Loadi #1071 to r[27]
  HD[812] = 32'b01100010101000000000000100000100;//Load m[#260] to r[21]
  HD[813] = 32'b01100110101000000000000011110001;//Store r[21] in m[#241]
  HD[814] = 32'b01010100000000000000001000010010;//Jump to #530
  HD[815] = 32'b01100010101000000000000011110010;//Load m[#242] to r[21]
  HD[816] = 32'b01100110101000000000000011101110;//Store r[21] in m[#238]
  HD[817] = 32'b01101011011000000000010000110011;//Loadi #1075 to r[27]
  HD[818] = 32'b01010100000000000000001000101110;//Jump to #558
  HD[819] = 32'b10001100000111000000000000000000;//Jump to r[28]
  HD[820] = 32'b01101100000000000000000000000000;//Nop
  HD[821] = 32'b01101100000000000000000000000000;//Nop
  HD[822] = 32'b01101100000000000000000000000000;//Nop
  HD[823] = 32'b01101100000000000000000000000000;//Nop
  HD[824] = 32'b01101100000000000000000000000000;//Nop
  HD[825] = 32'b01101100000000000000000000000000;//Nop
  HD[826] = 32'b01101100000000000000000000000000;//Nop
  HD[827] = 32'b01101011011000000000000100000001;//Loadi #257 to r[27]
  HD[828] = 32'b01010100000000000000010000111101;//Jump to #1085
  HD[829] = 32'b10100010101000000000000000000000;//Load wd to r[21]
  HD[830] = 32'b01100110101000000000000100001110;//Store r[21] in m[#270]
  HD[831] = 32'b01100010101000000000000100001110;//Load m[#270] to r[21]
  HD[832] = 32'b01011110110000001010100000000000;//SLT if r[0] < r[21], r[22] = 1 else r[22] = 0
  HD[833] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[834] = 32'b01001100000000000000000000001111;//Branch on Zero #15
  HD[835] = 32'b01101010111000000000000000000100;//Loadi #4 to r[23]
  HD[836] = 32'b01011110110101011011100000000000;//SLT if r[21] < r[23], r[22] = 1 else r[22] = 0
  HD[837] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[838] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[839] = 32'b01010100000000000000010001010100;//Jump to #1108
  HD[840] = 32'b01101010111000000000000000000101;//Loadi #5 to r[23]
  HD[841] = 32'b01011110110101011011100000000000;//SLT if r[21] < r[23], r[22] = 1 else r[22] = 0
  HD[842] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[843] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[844] = 32'b01010100000000000000010010111100;//Jump to #1212
  HD[845] = 32'b01101010111000000000000000000110;//Loadi #6 to r[23]
  HD[846] = 32'b01011110110101011011100000000000;//SLT if r[21] < r[23], r[22] = 1 else r[22] = 0
  HD[847] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[848] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[849] = 32'b01010100000000000000010100000100;//Jump to #1284
  HD[850] = 32'b01101100000000000000000000000000;//Nop
  HD[851] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[852] = 32'b01101100000000000000000000000000;//Nop
  HD[853] = 32'b01101100000000000000000000000000;//Nop
  HD[854] = 32'b01101100000000000000000000000000;//Nop
  HD[855] = 32'b01101100000000000000000000000000;//Nop
  HD[856] = 32'b01101100000000000000000000000000;//Nop
  HD[857] = 32'b01101011011000000000010010000011;//Loadi #1155 to r[27]
  HD[858] = 32'b01100010101000000000000100001110;//Load m[#270] to r[21]
  HD[859] = 32'b01100110101000000000000100010000;//Store r[21] in m[#272]
  HD[860] = 32'b01010100000000000000010001011101;//Jump to #1117
  HD[861] = 32'b01100100000000000000000100010010;//Store r[0] in m[#274]
  HD[862] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[863] = 32'b01100110101000000000000100010001;//Store r[21] in m[#273]
  HD[864] = 32'b01100010101000000000000100010001;//Load m[#273] to r[21]
  HD[865] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[866] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[867] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[868] = 32'b01001100000000000000000000011010;//Branch on Zero #26
  HD[869] = 32'b01101010111000000000000000000001;//Loadi #1 to r[23]
  HD[870] = 32'b01011110111101111011000000000000;//SLT if r[23] < r[22], r[23] = 1 else r[23] = 0
  HD[871] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[872] = 32'b01001100000000000000000000010011;//Branch on Zero #19
  HD[873] = 32'b00000110101101010000000000000011;//ADDi r[21], #3 to r[21]
  HD[874] = 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
  HD[875] = 32'b01011111000000001011100000000000;//SLT if r[0] < r[23], r[24] = 1 else r[24] = 0
  HD[876] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[877] = 32'b01001100000000000000000000001110;//Branch on Zero #14
  HD[878] = 32'b01101011000000000000000000000011;//Loadi #3 to r[24]
  HD[879] = 32'b01011111000101111100000000000000;//SLT if r[23] < r[24], r[24] = 1 else r[24] = 0
  HD[880] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[881] = 32'b01001100000000000000000000001010;//Branch on Zero #10
  HD[882] = 32'b00001110101101010000000000000010;//SUBi r[21], #2 to r[21]
  HD[883] = 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
  HD[884] = 32'b01100011000000000000000100010000;//Load m[#272] to r[24]
  HD[885] = 32'b01011110101101111100000000000000;//SLT if r[23] < r[24], r[21] = 1 else r[21] = 0
  HD[886] = 32'b01011111000110001011100000000000;//SLT if r[24] < r[23], r[24] = 1 else r[24] = 0
  HD[887] = 32'b00100111000101011100000000000000;//OR r[21],r[24] to r[24]
  HD[888] = 32'b00110111000110000000000000000000;//NOT r[24] to r[24]
  HD[889] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[890] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[891] = 32'b01100110110000000000000100010010;//Store r[22] in m[#274]
  HD[892] = 32'b01100010101000000000000100010001;//Load m[#273] to r[21]
  HD[893] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[894] = 32'b01010100000000000000010001011111;//Jump to #1119
  HD[895] = 32'b01101100000000000000000000000000;//Nop
  HD[896] = 32'b01101100000000000000000000000000;//Nop
  HD[897] = 32'b01101100000000000000000000000000;//Nop
  HD[898] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[899] = 32'b01101100000000000000000000000000;//Nop
  HD[900] = 32'b01101100000000000000000000000000;//Nop
  HD[901] = 32'b01100010101000000000000100010010;//Load m[#274] to r[21]
  HD[902] = 32'b01011110110000001010100000000000;//SLT if r[0] < r[21], r[22] = 1 else r[22] = 0
  HD[903] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[904] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[905] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[906] = 32'b10001100000111000000000000000000;//Jump to r[28]
  HD[907] = 32'b01101100000000000000000000000000;//Nop
  HD[908] = 32'b01101100000000000000000000000000;//Nop
  HD[909] = 32'b01101100000000000000000000000000;//Nop
  HD[910] = 32'b01100010101000000000000100010010;//Load m[#274] to r[21]
  HD[911] = 32'b01100110101000000000000100010011;//Store r[21] in m[#275]
  HD[912] = 32'b01101011011000000000010010101010;//Loadi #1194 to r[27]
  HD[913] = 32'b01010100000000000000010010010010;//Jump to #1170
  HD[914] = 32'b01100100000000000000000100010101;//Store r[0] in m[#277]
  HD[915] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[916] = 32'b01100110101000000000000100010100;//Store r[21] in m[#276]
  HD[917] = 32'b01100010101000000000000100010100;//Load m[#276] to r[21]
  HD[918] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[919] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[920] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[921] = 32'b01001100000000000000000000001101;//Branch on Zero #13
  HD[922] = 32'b01100010111000000000000100010011;//Load m[#275] to r[23]
  HD[923] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[924] = 32'b01011110111101111011000000000000;//SLT if r[23] < r[22], r[23] = 1 else r[23] = 0
  HD[925] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[926] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[927] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[928] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[929] = 32'b00000110101101010000000000000011;//ADDi r[21], #3 to r[21]
  HD[930] = 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
  HD[931] = 32'b01100110111000000000000100010101;//Store r[23] in m[#277]
  HD[932] = 32'b01100010101000000000000100010100;//Load m[#276] to r[21]
  HD[933] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[934] = 32'b01010100000000000000010010010100;//Jump to #1172
  HD[935] = 32'b01101100000000000000000000000000;//Nop
  HD[936] = 32'b01101100000000000000000000000000;//Nop
  HD[937] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[938] = 32'b01101100000000000000000000000000;//Nop
  HD[939] = 32'b01101100000000000000000000000000;//Nop
  HD[940] = 32'b01100010101000000000000100010101;//Load m[#277] to r[21]
  HD[941] = 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
  HD[942] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[943] = 32'b01011110110101101010100000000000;//SLT if r[22] < r[21], r[22] = 1 else r[22] = 0
  HD[944] = 32'b00100110110101101011100000000000;//OR r[22],r[23] to r[22]
  HD[945] = 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
  HD[946] = 32'b01111100000101100000000000000000;//Pre Branch r[22]
  HD[947] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[948] = 32'b10001100000111000000000000000000;//Jump to r[28]
  HD[949] = 32'b01100010101000000000000100010010;//Load m[#274] to r[21]
  HD[950] = 32'b01100110101000000000000100000101;//Store r[21] in m[#261]
  HD[951] = 32'b01100110101000000000000100000100;//Store r[21] in m[#260]
  HD[952] = 32'b01101011011000000000001111001101;//Loadi #973 to r[27]
  HD[953] = 32'b01010100000000000000001110101101;//Jump to #941
  HD[954] = 32'b01101100000000000000000000000000;//Nop
  HD[955] = 32'b01101100000000000000000000000000;//Nop
  HD[956] = 32'b01101100000000000000000000000000;//Nop
  HD[957] = 32'b01101100000000000000000000000000;//Nop
  HD[958] = 32'b01101011011000000000010011000000;//Loadi #1216 to r[27]
  HD[959] = 32'b01010100000000000000001010000011;//Jump to #643
  HD[960] = 32'b01100010101000000000000100001111;//Load m[#271] to r[21]
  HD[961] = 32'b01100010110000000000000011110111;//Load m[#247] to r[22]
  HD[962] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[963] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[964] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[965] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[966] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[967] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[968] = 32'b00000111100111000000000000000001;//ADDi r[28], #1 to r[28]
  HD[969] = 32'b10001100000111000000000000000000;//Jump to r[28]
  HD[970] = 32'b01101100000000000000000000000000;//Nop
  HD[971] = 32'b01101100000000000000000000000000;//Nop
  HD[972] = 32'b00000111100111000000000000000001;//ADDi r[28], #1 to r[28]
  HD[973] = 32'b01101011011000000000010011010110;//Loadi #1238 to r[27]
  HD[974] = 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
  HD[975] = 32'b01100110101000000000000011100100;//Store r[21] in m[#228]
  HD[976] = 32'b01100100000000000000000011100101;//Store r[0] in m[#229]
  HD[977] = 32'b01100100000000000000000011100110;//Store r[0] in m[#230]
  HD[978] = 32'b01101010101000000000000000000010;//Loadi #2 to r[21]
  HD[979] = 32'b01100110101000000000000011100111;//Store r[21] in m[#231]
  HD[980] = 32'b01100111100000000000000011101000;//Store r[28] in m[#232]
  HD[981] = 32'b01010100000000000000000111001101;//Jump to #461
  HD[982] = 32'b01101100000000000000000000000000;//Nop
  HD[983] = 32'b01101100000000000000000000000000;//Nop
  HD[984] = 32'b01100010101000000000000100001111;//Load m[#271] to r[21]
  HD[985] = 32'b01100110101000000000000100000101;//Store r[21] in m[#261]
  HD[986] = 32'b01100110101000000000000100000100;//Store r[21] in m[#260]
  HD[987] = 32'b01101011011000000000001111001101;//Loadi #973 to r[27]
  HD[988] = 32'b01010100000000000000001110101101;//Jump to #941
  HD[989] = 32'b01101100000000000000000000000000;//Nop
  HD[990] = 32'b01101100000000000000000000000000;//Nop
  HD[991] = 32'b01101100000000000000000000000000;//Nop
  HD[992] = 32'b01101100000000000000000000000000;//Nop
  HD[993] = 32'b01100110101000000000000100010111;//Store r[21] in m[#279]
  HD[994] = 32'b01101010110000000000000000000100;//Loadi #4 to r[22]
  HD[995] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[996] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[997] = 32'b01001100000000000000000000011010;//Branch on Zero #26
  HD[998] = 32'b01101011011000000000010011111101;//Loadi #1277 to r[27]
  HD[999] = 32'b01010100000000000000010011101000;//Jump to #1256
  HD[1000] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[1001] = 32'b01100110101000000000000100010110;//Store r[21] in m[#278]
  HD[1002] = 32'b01100010101000000000000100010110;//Load m[#278] to r[21]
  HD[1003] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[1004] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[1005] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[1006] = 32'b01001100000000000000000000001011;//Branch on Zero #11
  HD[1007] = 32'b00000110101101010000000000000011;//ADDi r[21], #3 to r[21]
  HD[1008] = 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
  HD[1009] = 32'b01101010101000000000000000000010;//Loadi #2 to r[21]
  HD[1010] = 32'b01011111000101111010100000000000;//SLT if r[23] < r[21], r[24] = 1 else r[24] = 0
  HD[1011] = 32'b00110111000110000000000000000000;//NOT r[24] to r[24]
  HD[1012] = 32'b01111100000110000000000000000000;//Pre Branch r[24]
  HD[1013] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[1014] = 32'b10000010110000000000000000000000;//Output r[22]
  HD[1015] = 32'b01100010101000000000000100010110;//Load m[#278] to r[21]
  HD[1016] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[1017] = 32'b01010100000000000000010011101001;//Jump to #1257
  HD[1018] = 32'b01101100000000000000000000000000;//Nop
  HD[1019] = 32'b01101100000000000000000000000000;//Nop
  HD[1020] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[1021] = 32'b01101100000000000000000000000000;//Nop
  HD[1022] = 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
  HD[1023] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[1024] = 32'b01101100000000000000000000000000;//Nop
  HD[1025] = 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
  HD[1026] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[1027] = 32'b01101100000000000000000000000000;//Nop
  HD[1028] = 32'b01101100000000000000000000000000;//Nop
  HD[1029] = 32'b01101100000000000000000000000000;//Nop
  HD[1030] = 32'b01101100000000000000000000000000;//Nop
  HD[1031] = 32'b01101100000000000000000000000000;//Nop
  HD[1032] = 32'b01101011011000000000010100001010;//Loadi #1290 to r[27]
  HD[1033] = 32'b01010100000000000000001010000011;//Jump to #643
  HD[1034] = 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
  HD[1035] = 32'b01100110101000000000000011100100;//Store r[21] in m[#228]
  HD[1036] = 32'b01100100000000000000000011100101;//Store r[0] in m[#229]
  HD[1037] = 32'b01100100000000000000000011100110;//Store r[0] in m[#230]
  HD[1038] = 32'b01100100000000000000000011100111;//Store r[0] in m[#231]
  HD[1039] = 32'b01100100000000000000000011101000;//Store r[0] in m[#232]
  HD[1040] = 32'b01101011011000000000010100010010;//Loadi #1298 to r[27]
  HD[1041] = 32'b01010100000000000000000111001101;//Jump to #461
  HD[1042] = 32'b01101100000000000000000000000000;//Nop
  HD[1043] = 32'b01101100000000000000000000000000;//Nop
  HD[1044] = 32'b01101100000000000000000000000000;//Nop
  HD[1045] = 32'b01101100000000000000000000000000;//Nop
  HD[1046] = 32'b01101011011000000000010100110000;//Loadi #1328 to r[27]
  HD[1047] = 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
  HD[1048] = 32'b01100110101000000000000100011000;//Store r[21] in m[#280]
  HD[1049] = 32'b01010100000000000000010100011010;//Jump to #1306
  HD[1050] = 32'b01101010101000000000000011000000;//Loadi #192 to r[21]
  HD[1051] = 32'b01100110101000000000000100011001;//Store r[21] in m[#281]
  HD[1052] = 32'b01100010101000000000000100011001;//Load m[#281] to r[21]
  HD[1053] = 32'b10000110110101010000000000000000;//Loadr m[r[21]] to r[22]
  HD[1054] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[1055] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[1056] = 32'b01001100000000000000000000001100;//Branch on Zero #12
  HD[1057] = 32'b01100010111000000000000100011000;//Load m[#280] to r[23]
  HD[1058] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[1059] = 32'b01011110111101111011000000000000;//SLT if r[23] < r[22], r[23] = 1 else r[23] = 0
  HD[1060] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[1061] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[1062] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[1063] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[1064] = 32'b01101010111000000000000000000001;//Loadi #1 to r[23]
  HD[1065] = 32'b10001010111101010000000000000000;//rStore r[23] in m[r[21]]
  HD[1066] = 32'b01100010101000000000000100011001;//Load m[#281] to r[21]
  HD[1067] = 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
  HD[1068] = 32'b01010100000000000000010100011011;//Jump to #1307
  HD[1069] = 32'b01101100000000000000000000000000;//Nop
  HD[1070] = 32'b01101100000000000000000000000000;//Nop
  HD[1071] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[1072] = 32'b01101100000000000000000000000000;//Nop
  HD[1073] = 32'b01101100000000000000000000000000;//Nop
  HD[1074] = 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
  HD[1075] = 32'b01100010110000000000000100001111;//Load m[#271] to r[22]
  HD[1076] = 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
  HD[1077] = 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
  HD[1078] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[1079] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[1080] = 32'b01001100000000000000000000001000;//Branch on Zero #8
  HD[1081] = 32'b01100010101000000000000100001111;//Load m[#271] to r[21]
  HD[1082] = 32'b01100110101000000000000100000101;//Store r[21] in m[#261]
  HD[1083] = 32'b01100110101000000000000100000100;//Store r[21] in m[#260]
  HD[1084] = 32'b01101011011000000000001111001101;//Loadi #973 to r[27]
  HD[1085] = 32'b01010100000000000000001110101101;//Jump to #941
  HD[1086] = 32'b01101100000000000000000000000000;//Nop
  HD[1087] = 32'b01101100000000000000000000000000;//Nop
  HD[1088] = 32'b01101100000000000000000000000000;//Nop
  HD[1089] = 32'b01010100000000000000000100000000;//Jump to #256
  HD[1090] = 32'b01101100000000000000000000000000;//Nop
  HD[1091] = 32'b01100010110000000000000100000111;//Load m[#263] to r[22]
  HD[1092] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[1093] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[1094] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[1095] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[1096] = 32'b10001100000111000000000000000000;//Jump to r[28]
  HD[1097] = 32'b01010100000000000000001111001101;//Jump to #973
  HD[1098] = 32'b01101100000000000000000000000000;//Nop
  HD[1099] = 32'b01101100000000000000000000000000;//Nop
  HD[1100] = 32'b01100010101000000000000100000100;//Load m[#260] to r[21]
  HD[1101] = 32'b01100110101000000000000011100100;//Store r[21] in m[#228]
  HD[1102] = 32'b01100100000000000000000011100101;//Store r[0] in m[#229]
  HD[1103] = 32'b01100100000000000000000011100110;//Store r[0] in m[#230]
  HD[1104] = 32'b01100100000000000000000011100111;//Store r[0] in m[#231]
  HD[1105] = 32'b01100100000000000000000011101000;//Store r[0] in m[#232]
  HD[1106] = 32'b01101011011000000000010101010101;//Loadi #1365 to r[27]
  HD[1107] = 32'b01010100000000000000000111001101;//Jump to #461
  HD[1108] = 32'b01101100000000000000000000000000;//Nop
  HD[1109] = 32'b01101100000000000000000000000000;//Nop
  HD[1110] = 32'b01101100000000000000000000000000;//Nop
  HD[1111] = 32'b01100010101000000000000100000100;//Load m[#260] to r[21]
  HD[1112] = 32'b01100110101000000000000100011000;//Store r[21] in m[#280]
  HD[1113] = 32'b01101011011000000000010101011011;//Loadi #1371 to r[27]
  HD[1114] = 32'b01010100000000000000010100011010;//Jump to #1306
  HD[1115] = 32'b01010100000000000000000100000001;//Jump to #257
  HD[1116] = 32'b01101100000000000000000000000000;//Nop
  HD[1117] = 32'b01101100000000000000000000000000;//Nop
  HD[1118] = 32'b01101100000000000000000000000000;//Nop
  HD[1119] = 32'b01110110101000000000000000000000;//Input to r[21]
  HD[1120] = 32'b01100110101000000000000100011011;//Store r[21] in m[#283]
  HD[1121] = 32'b01100010101000000000000011101010;//Load m[#234] to r[21]
  HD[1122] = 32'b01100110101000000000000100011010;//Store r[21] in m[#282]
  HD[1123] = 32'b01101011011000000000010101111100;//Loadi #1404 to r[27]
  HD[1124] = 32'b01010100000000000000010101100101;//Jump to #1381
  HD[1125] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[1126] = 32'b01101010101000000000100000000000;//Loadi #1, #0 to r[21]
  HD[1127] = 32'b01100110101000000000000100011100;//Store r[21] in m[#284]
  HD[1128] = 32'b01100010101000000000000100011100;//Load m[#284] to r[21]
  HD[1129] = 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
  HD[1130] = 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
  HD[1131] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[1132] = 32'b01001100000000000000000000001100;//Branch on Zero #12
  HD[1133] = 32'b01100010111000000000000100011010;//Load m[#282] to r[23]
  HD[1134] = 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
  HD[1135] = 32'b01011110111101111011000000000000;//SLT if r[23] < r[22], r[23] = 1 else r[23] = 0
  HD[1136] = 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
  HD[1137] = 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
  HD[1138] = 32'b01111100000101110000000000000000;//Pre Branch r[23]
  HD[1139] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[1140] = 32'b01100010111000000000000100011011;//Load m[#283] to r[23]
  HD[1141] = 32'b10010010111101010000000000000000;//hdStore r[23] in m[r[21]]
  HD[1142] = 32'b01010100000000000000010101111001;//Jump to #1401
  HD[1143] = 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
  HD[1144] = 32'b01010100000000000000010101100111;//Jump to #1383
  HD[1145] = 32'b01101100000000000000000000000000;//Nop
  HD[1146] = 32'b01101100000000000000000000000000;//Nop
  HD[1147] = 32'b10001100000110110000000000000000;//Jump to r[27]
  HD[1148] = 32'b01101100000000000000000000000000;//Nop
  HD[1149] = 32'b01010100000000000000000100101011;//Jump to #299
  HD[1150] = 32'b01110000000000000000000000000000;//Hlt
  HD[1151] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]




//programs & processess' list of information
//program 0 [line 2048]
		 HD[2048] = 32'b00000000000000000000000000001011;
     HD[2049] = 32'b00000000000000000000000000000000;
     HD[2051] = 32'b00000000000000000000000000000000;
     HD[2053] = 32'b00000000000000000000000000000000;

//program 1 [line 2080]
		 HD[2080] = 32'b00000000000000000000000000001100;
		 HD[2081] = 32'b00000000000000000000000000000000;
     HD[2083] = 32'b00000000000000000000000000000000;
		 HD[2085] = 32'b00000000000000000000000000000001;

//program 2 [line 2112]
		 HD[2112] = 32'b00000000000000000000000000001101;
		 HD[2113] = 32'b00000000000000000000000000000000;
		 HD[2115] = 32'b00000000000000000000000000000000;
		 HD[2117] = 32'b00000000000000000000000000000010;

//program 3 [line 2144]
		 HD[2144] = 32'b00000000000000000000000000001110;
		 HD[2145] = 32'b00000000000000000000000000000000;
		 HD[2147] = 32'b00000000000000000000000000000000;
		 HD[2149] = 32'b00000000000000000000000000000011;

//program 4 [line 2176]
		 HD[2176] = 32'b00000000000000000000000000001111;
		 HD[2177] = 32'b00000000000000000000000000000000;
		 HD[2179] = 32'b00000000000000000000000000000000;
     HD[2181] = 32'b00000000000000000000000000000100;

 //program 5 [line 2208]
     HD[2208] = 32'b00000000000000000000000000010000;
     HD[2209] = 32'b00000000000000000000000000000000;
     HD[2211] = 32'b00000000000000000000000000000000;
     HD[2213] = 32'b00000000000000000000000000000101;

 //program 6 [line 2240]
     HD[2240] = 32'b00000000000000000000000000010001;
     HD[2241] = 32'b00000000000000000000000000000000;
     HD[2243] = 32'b00000000000000000000000000000000;
     HD[2245] = 32'b00000000000000000000000000000110;

 //program 7 [line 2272]
     HD[2272] = 32'b00000000000000000000000000010010;
     HD[2273] = 32'b00000000000000000000000000000000;
     HD[2275] = 32'b00000000000000000000000000000000;
     HD[2277] = 32'b00000000000000000000000000000111;

 //program 8 [line 2304]
     HD[2304] = 32'b00000000000000000000000000010011;
     HD[2305] = 32'b00000000000000000000000000000000;
     HD[2307] = 32'b00000000000000000000000000000000;
     HD[2309] = 32'b00000000000000000000000000001000;

 //program 9 [line 2336]
     HD[2336] = 32'b00000000000000000000000000010100;
     HD[2337] = 32'b00000000000000000000000000000000;
     HD[2339] = 32'b00000000000000000000000000000000;
     HD[2341] = 32'b00000000000000000000000000001001;


//programs' instructions
//program 0 [line 4096] - Fibonacci
HD[4096] = 32'b01101100000000000000000000000000;//Nop
HD[4097] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
HD[4098] = 32'b01111000000000000000000000000000;//preio
HD[4099] = 32'b01110100001000000000000000000000;//Input to r[1]
HD[4100] = 32'b01100100001000000000000000000010;//Store r[1] in m[#2]
HD[4101] = 32'b01100100000000000000000000000101;//Store r[0] in m[#5]
HD[4102] = 32'b01101000001000000000000000000001;//Loadi #1 to r[1]
HD[4103] = 32'b01100100001000000000000000000110;//Store r[1] in m[#6]
HD[4104] = 32'b01100100000000000000000000000011;//Store r[0] in m[#3]
HD[4105] = 32'b01100000001000000000000000000010;//Load m[#2] to r[1]
HD[4106] = 32'b00000100001000010000000000000001;//ADDi r[1], #1 to r[1]
HD[4107] = 32'b01100000010000000000000000000011;//Load m[#3] to r[2]
HD[4108] = 32'b01100100010000000000000000000011;//Store r[2] in m[#3]
HD[4109] = 32'b01011100100000100000100000000000;//SLT if r[2] < r[1], r[4] = 1 else r[4] = 0
HD[4110] = 32'b01111100000001000000000000000000;//Pre Branch r[4]
HD[4111] = 32'b01001100000000000000000000010000;//Branch on Zero #16
HD[4112] = 32'b01101000110000000000000000000010;//Loadi #2 to r[6]
HD[4113] = 32'b01011100100000100011000000000000;//SLT if r[2] < r[6], r[4] = 1 else r[4] = 0
HD[4114] = 32'b01111100000001000000000000000000;//Pre Branch r[4]
HD[4115] = 32'b01001100000000000000000000000011;//Branch on Zero #3
HD[4116] = 32'b01100001000000000000000000000011;//Load m[#3] to r[8]
HD[4117] = 32'b01100101000000000000000000000100;//Store r[8] in m[#4]
HD[4118] = 32'b01010100000000000000000000011101;//Jump to #29
HD[4119] = 32'b01100001000000000000000000000101;//Load m[#5] to r[8]
HD[4120] = 32'b01100001001000000000000000000110;//Load m[#6] to r[9]
HD[4121] = 32'b00000001000010000100100000000000;//ADD r[8],r[9] to r[8]
HD[4122] = 32'b01100101000000000000000000000100;//Store r[8] in m[#4]
HD[4123] = 32'b01100101001000000000000000000101;//Store r[9] in m[#5]
HD[4124] = 32'b01100101000000000000000000000110;//Store r[8] in m[#6]
HD[4125] = 32'b01100000010000000000000000000011;//Load m[#3] to r[2]
HD[4126] = 32'b00000100010000100000000000000001;//ADDi r[2], #1 to r[2]
HD[4127] = 32'b01010100000000000000000000001100;//Jump to #12
HD[4128] = 32'b01100000101000000000000000000100;//Load m[#4] to r[5]
HD[4129] = 32'b01111000000000000000000000000000;//preio
HD[4130] = 32'b10000000101000000000000000000000;//Output r[5]
HD[4131] = 32'b01110000000000000000000000000000;//Hlt
HD[4132] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]




//program 1 [line 4288] - Biggest
	 	 HD[4288] = 32'b01101100000000000000000000000000;//Nop
	 	 HD[4289] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
	 	 HD[4290] = 32'b01101001011000000000000000000011;//Loadi #3 to r[11]
	 	 HD[4291] = 32'b01100101011000000000000000000100;//Store r[11] in m[#4]
	 	 HD[4292] = 32'b01100100000000000000000000000101;//Store r[0] in m[#5]
	 	 HD[4293] = 32'b01111000000000000000000000000000;//preio
	 	 HD[4294] = 32'b01110101011000000000000000000000;//Input to r[11]
	 	 HD[4295] = 32'b01100101011000000000000000000001;//Store r[11] in m[#1]
	 	 HD[4296] = 32'b01111000000000000000000000000000;//preio
	 	 HD[4297] = 32'b01110101011000000000000000000000;//Input to r[11]
	 	 HD[4298] = 32'b01100101011000000000000000000010;//Store r[11] in m[#2]
	 	 HD[4299] = 32'b01111000000000000000000000000000;//preio
	 	 HD[4300] = 32'b01110101011000000000000000000000;//Input to r[11]
	 	 HD[4301] = 32'b01100101011000000000000000000011;//Store r[11] in m[#3]
	 	 HD[4302] = 32'b01100100000000000000000000000110;//Store r[0] in m[#6]
	 	 HD[4303] = 32'b01100100000000000000000000000111;//Store r[0] in m[#7]
	 	 HD[4304] = 32'b01100001100000000000000000000100;//Load m[#4] to r[12]
	 	 HD[4305] = 32'b01100001011000000000000000000111;//Load m[#7] to r[11]
	 	 HD[4306] = 32'b01011101101010110110000000000000;//SLT if r[11] < r[12], r[13] = 1 else r[13] = 0
	 	 HD[4307] = 32'b01111100000011010000000000000000;//Pre Branch r[13]
	 	 HD[4308] = 32'b01001100000000000000000000001010;//Branch on Zero #10
	 	 HD[4309] = 32'b01100001101000000000000000000110;//Load m[#6] to r[13]
	 	 HD[4310] = 32'b00000101110010110000000000000001;//ADDi r[11], #1 to r[14]
	 	 HD[4311] = 32'b10000101110011100000000000000000;//Loadr m[r[14]] to r[14]
	 	 HD[4312] = 32'b01011101111011010111000000000000;//SLT if r[13] < r[14], r[15] = 1 else r[15] = 0
	 	 HD[4313] = 32'b01111100000011110000000000000000;//Pre Branch r[15]
	 	 HD[4314] = 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[4315] = 32'b01100101110000000000000000000110;//Store r[14] in m[#6]
	 	 HD[4316] = 32'b00000101011010110000000000000001;//ADDi r[11], #1 to r[11]
	 	 HD[4317] = 32'b01100101011000000000000000000111;//Store r[11] in m[#7]
	 	 HD[4318] = 32'b01010100000000000000000000010001;//Jump to #17
	 	 HD[4319] = 32'b01100000101000000000000000000110;//Load m[#6] to r[5]
	 	 HD[4320] = 32'b01111000000000000000000000000000;//preio
	 	 HD[4321] = 32'b10000000101000000000000000000000;//Output r[5]
	 	 HD[4322] = 32'b01110000000000000000000000000000;//Hlt
	 	 HD[4323] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]





//program 2 [line 4480] - Division [13]
HD[4480] = 32'b01101100000000000000000000000000;//Nop
HD[4481] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
HD[4482] = 32'b01100100000000000000000000000011;//Store r[0] in m[#3]
HD[4483] = 32'b01111000000000000000000000000000;//preio
HD[4484] = 32'b01110101011000000000000000000000;//Input to r[11]
HD[4485] = 32'b01100101011000000000000000000001;//Store r[11] in m[#1]
HD[4486] = 32'b01111000000000000000000000000000;//preio
HD[4487] = 32'b01110101011000000000000000000000;//Input to r[11]
HD[4488] = 32'b01100101011000000000000000000010;//Store r[11] in m[#2]
HD[4489] = 32'b01100001011000000000000000000001;//Load m[#1] to r[11]
HD[4490] = 32'b01100001100000000000000000000010;//Load m[#2] to r[12]
HD[4491] = 32'b00000101111010110000000000000001;//ADDi r[11], #1 to r[15]
HD[4492] = 32'b01011101111011000111100000000000;//SLT if r[12] < r[15], r[15] = 1 else r[15] = 0
HD[4493] = 32'b01111100000011110000000000000000;//Pre Branch r[15]
HD[4494] = 32'b01001100000000000000000000000110;//Branch on Zero #6
HD[4495] = 32'b00001001011010110110000000000000;//SUB r[11],r[12] to r[11]
HD[4496] = 32'b01100101011000000000000000000001;//Store r[11] in m[#1]
HD[4497] = 32'b01100001101000000000000000000011;//Load m[#3] to r[13]
HD[4498] = 32'b00000101101011010000000000000001;//ADDi r[13], #1 to r[13]
HD[4499] = 32'b01100101101000000000000000000011;//Store r[13] in m[#3]
HD[4500] = 32'b01010100000000000000000000001001;//Jump to #9
HD[4501] = 32'b01100001101000000000000000000011;//Load m[#3] to r[13]
HD[4502] = 32'b01111000000000000000000000000000;//preio
HD[4503] = 32'b10000001101000000000000000000000;//Output r[13]
HD[4504] = 32'b01110000000000000000000000000000;//Hlt
HD[4505] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]



  //program 3 [line 4672] - Pow [14]
  HD[4672] = 32'b01101100000000000000000000000000;//Nop
  HD[4673] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[4674] = 32'b01111000000000000000000000000000;//preio
  HD[4675] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[4676] = 32'b01100101011000000000000000000010;//Store r[11] in m[#2]
  HD[4677] = 32'b01111000000000000000000000000000;//preio
  HD[4678] = 32'b01110101100000000000000000000000;//Input to r[12]
  HD[4679] = 32'b01100101100000000000000000000011;//Store r[12] in m[#3]
  HD[4680] = 32'b01101001101000000000000000000001;//Loadi #1 to r[13]
  HD[4681] = 32'b01100101101000000000000000000100;//Store r[13] in m[#4]
  HD[4682] = 32'b01100001011000000000000000000011;//Load m[#3] to r[11]
  HD[4683] = 32'b01011101100000000101100000000000;//SLT if r[0] < r[11], r[12] = 1 else r[12] = 0
  HD[4684] = 32'b01111100000011000000000000000000;//Pre Branch r[12]
  HD[4685] = 32'b01001100000000000000000000000110;//Branch on Zero #6
  HD[4686] = 32'b01100001110000000000000000000100;//Load m[#4] to r[14]
  HD[4687] = 32'b01100001100000000000000000000010;//Load m[#2] to r[12]
  HD[4688] = 32'b00010001111011000111000000000000;//TIMES r[12],r[14] to r[15]
  HD[4689] = 32'b01100101111000000000000000000100;//Store r[15] in m[#4]
  HD[4690] = 32'b00001101011010110000000000000001;//SUBi r[11], #1 to r[11]
  HD[4691] = 32'b01010100000000000000000000001011;//Jump to #11
  HD[4692] = 32'b01100001000000000000000000000100;//Load m[#4] to r[8]
  HD[4693] = 32'b01111000000000000000000000000000;//preio
  HD[4694] = 32'b10000001000000000000000000000000;//Output r[8]
  HD[4695] = 32'b01110000000000000000000000000000;//Hlt
  HD[4696] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]




  //program 4 [line 4864] - Mean [15]
  HD[4864] = 32'b01101100000000000000000000000000;//Nop
  HD[4865] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[4866] = 32'b01111000000000000000000000000000;//preio
  HD[4867] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[4868] = 32'b01100101011000000000000000000010;//Store r[11] in m[#2]
  HD[4869] = 32'b01111000000000000000000000000000;//preio
  HD[4870] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[4871] = 32'b01100101011000000000000000000011;//Store r[11] in m[#3]
  HD[4872] = 32'b01111000000000000000000000000000;//preio
  HD[4873] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[4874] = 32'b01100101011000000000000000000100;//Store r[11] in m[#4]
  HD[4875] = 32'b01100100000000000000000000000111;//Store r[0] in m[#7]
  HD[4876] = 32'b01100100000000000000000000000110;//Store r[0] in m[#6]
  HD[4877] = 32'b01101001011000000000000000000011;//Loadi #3 to r[11]
  HD[4878] = 32'b01100101011000000000000000000101;//Store r[11] in m[#5]
  HD[4879] = 32'b01100001100000000000000000000110;//Load m[#6] to r[12]
  HD[4880] = 32'b01100001010000000000000000000101;//Load m[#5] to r[10]
  HD[4881] = 32'b01011101101011000101000000000000;//SLT if r[12] < r[10], r[13] = 1 else r[13] = 0
  HD[4882] = 32'b01111100000011010000000000000000;//Pre Branch r[13]
  HD[4883] = 32'b01001100000000000000000000000111;//Branch on Zero #7
  HD[4884] = 32'b00000100010011000000000000000010;//ADDi r[12], #2 to r[2]
  HD[4885] = 32'b10000100010000100000000000000000;//Loadr m[r[2]] to r[2]
  HD[4886] = 32'b01100001110000000000000000000111;//Load m[#7] to r[14]
  HD[4887] = 32'b00000000010000100111000000000000;//ADD r[2],r[14] to r[2]
  HD[4888] = 32'b01100100010000000000000000000111;//Store r[2] in m[#7]
  HD[4889] = 32'b00000101100011000000000000000001;//ADDi r[12], #1 to r[12]
  HD[4890] = 32'b01010100000000000000000000010001;//Jump to #17
  HD[4891] = 32'b01100001110000000000000000000111;//Load m[#7] to r[14]
  HD[4892] = 32'b01100001010000000000000000000101;//Load m[#5] to r[10]
  HD[4893] = 32'b00010101101011100101000000000000;//DIVIDE r[14],r[10] to r[13]
  HD[4894] = 32'b01111000000000000000000000000000;//preio
  HD[4895] = 32'b10000001101000000000000000000000;//Output r[13]
  HD[4896] = 32'b01110000000000000000000000000000;//Hlt
  HD[4897] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]



  //program 5 [line 5056] - Smallest [16]
  HD[5056] = 32'b01101100000000000000000000000000;//Nop
  HD[5057] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[5058] = 32'b01101001011000000000000000000011;//Loadi #3 to r[11]
  HD[5059] = 32'b01100101011000000000000000000100;//Store r[11] in m[#4]
  HD[5060] = 32'b01100100000000000000000000000101;//Store r[0] in m[#5]
  HD[5061] = 32'b01111000000000000000000000000000;//preio
  HD[5062] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[5063] = 32'b01100101011000000000000000000001;//Store r[11] in m[#1]
  HD[5064] = 32'b01111000000000000000000000000000;//preio
  HD[5065] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[5066] = 32'b01100101011000000000000000000010;//Store r[11] in m[#2]
  HD[5067] = 32'b01111000000000000000000000000000;//preio
  HD[5068] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[5069] = 32'b01100101011000000000000000000011;//Store r[11] in m[#3]
  HD[5070] = 32'b01101001011000111101000010010000;//Loadi #250000 to r[11]
  HD[5071] = 32'b01100101011000000000000000000110;//Store r[11] in m[#6]
  HD[5072] = 32'b01100100000000000000000000000111;//Store r[0] in m[#7]
  HD[5073] = 32'b01100001100000000000000000000100;//Load m[#4] to r[12]
  HD[5074] = 32'b01100001011000000000000000000111;//Load m[#7] to r[11]
  HD[5075] = 32'b01011101101010110110000000000000;//SLT if r[11] < r[12], r[13] = 1 else r[13] = 0
  HD[5076] = 32'b01111100000011010000000000000000;//Pre Branch r[13]
  HD[5077] = 32'b01001100000000000000000000001011;//Branch on Zero #11
  HD[5078] = 32'b01100001101000000000000000000110;//Load m[#6] to r[13]
  HD[5079] = 32'b00000101110010110000000000000001;//ADDi r[11], #1 to r[14]
  HD[5080] = 32'b10000101110011100000000000000000;//Loadr m[r[14]] to r[14]
  HD[5081] = 32'b01011101111011100110100000000000;//SLT if r[14] < r[13], r[15] = 1 else r[15] = 0
  HD[5082] = 32'b01111100000011110000000000000000;//Pre Branch r[15]
  HD[5083] = 32'b01001100000000000000000000000001;//Branch on Zero #1
  HD[5084] = 32'b01100101110000000000000000000110;//Store r[14] in m[#6]
  HD[5085] = 32'b00000101011010110000000000000001;//ADDi r[11], #1 to r[11]
  HD[5086] = 32'b01101100000000000000000000000000;//Nop
  HD[5087] = 32'b01100101011000000000000000000111;//Store r[11] in m[#7]
  HD[5088] = 32'b01010100000000000000000000010010;//Jump to #18
  HD[5089] = 32'b01100000101000000000000000000110;//Load m[#6] to r[5]
  HD[5090] = 32'b01111000000000000000000000000000;//preio
  HD[5091] = 32'b10000000101000000000000000000000;//Output r[5]
  HD[5092] = 32'b01110000000000000000000000000000;//Hlt
  HD[5093] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]


  //program 6 [line 5248] - Sort [17]
  HD[5248] = 32'b01101100000000000000000000000000;//Nop
  HD[5249] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[5250] = 32'b01111000000000000000000000000000;//preio
  HD[5251] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[5252] = 32'b01100101011000000000000000000000;//Store r[11] in m[#0]
  HD[5253] = 32'b01111000000000000000000000000000;//preio
  HD[5254] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[5255] = 32'b01100101011000000000000000000001;//Store r[11] in m[#1]
  HD[5256] = 32'b01111000000000000000000000000000;//preio
  HD[5257] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[5258] = 32'b01100101011000000000000000000010;//Store r[11] in m[#2]
  HD[5259] = 32'b01111000000000000000000000000000;//preio
  HD[5260] = 32'b01110101011000000000000000000000;//Input to r[11]
  HD[5261] = 32'b01100101011000000000000000000011;//Store r[11] in m[#3]
  HD[5262] = 32'b01100100000000000000000000000100;//Store r[0] in m[#4]
  HD[5263] = 32'b01101001011000000000000000000100;//Loadi #4 to r[11]
  HD[5264] = 32'b01100101011000000000000000001000;//Store r[11] in m[#8]
  HD[5265] = 32'b01100001000000000000000000000100;//Load m[#4] to r[8]
  HD[5266] = 32'b01100010000000000000000000001000;//Load m[#8] to r[16]
  HD[5267] = 32'b00001101111100000000000000000001;//SUBi r[16], #1 to r[15]
  HD[5268] = 32'b01011101111010000111100000000000;//SLT if r[8] < r[15], r[15] = 1 else r[15] = 0
  HD[5269] = 32'b01111100000011110000000000000000;//Pre Branch r[15]
  HD[5270] = 32'b01001100000000000000000000100110;//Branch on Zero #38
  HD[5271] = 32'b01100101000000000000000000000110;//Store r[8] in m[#6]
  HD[5272] = 32'b00000001001010000000000000000000;//ADD r[8],r[0] to r[9]
  HD[5273] = 32'b01100101001000000000000000000101;//Store r[9] in m[#5]
  HD[5274] = 32'b01100001010000000000000000000101;//Load m[#5] to r[10]
  HD[5275] = 32'b01011101111010101000000000000000;//SLT if r[10] < r[16], r[15] = 1 else r[15] = 0
  HD[5276] = 32'b01111100000011110000000000000000;//Pre Branch r[15]
  HD[5277] = 32'b01001100000000000000000000001100;//Branch on Zero #12
  HD[5278] = 32'b01100001100000000000000000000110;//Load m[#6] to r[12]
  HD[5279] = 32'b10000101010010100000000000000000;//Loadr m[r[10]] to r[10]
  HD[5280] = 32'b10000101100011000000000000000000;//Loadr m[r[12]] to r[12]
  HD[5281] = 32'b01011101011010100110000000000000;//SLT if r[10] < r[12], r[11] = 1 else r[11] = 0
  HD[5282] = 32'b01111100000010110000000000000000;//Pre Branch r[11]
  HD[5283] = 32'b01001100000000000000000000000010;//Branch on Zero #2
  HD[5284] = 32'b01100001010000000000000000000101;//Load m[#5] to r[10]
  HD[5285] = 32'b01100101010000000000000000000110;//Store r[10] in m[#6]
  HD[5286] = 32'b01100001010000000000000000000101;//Load m[#5] to r[10]
  HD[5287] = 32'b00000101010010100000000000000001;//ADDi r[10], #1 to r[10]
  HD[5288] = 32'b01100101010000000000000000000101;//Store r[10] in m[#5]
  HD[5289] = 32'b01010100000000000000000000011010;//Jump to #26
  HD[5290] = 32'b01100001000000000000000000000100;//Load m[#4] to r[8]
  HD[5291] = 32'b01100001100000000000000000000110;//Load m[#6] to r[12]
  HD[5292] = 32'b01011101011010000110000000000000;//SLT if r[8] < r[12], r[11] = 1 else r[11] = 0
  HD[5293] = 32'b01011101101011000100000000000000;//SLT if r[12] < r[8], r[13] = 1 else r[13] = 0
  HD[5294] = 32'b00100101011010110110100000000000;//OR r[11],r[13] to r[11]
  HD[5295] = 32'b01111100000010110000000000000000;//Pre Branch r[11]
  HD[5296] = 32'b01001100000000000000000000001000;//Branch on Zero #8
  HD[5297] = 32'b10000101000010000000000000000000;//Loadr m[r[8]] to r[8]
  HD[5298] = 32'b01100101000000000000000000000111;//Store r[8] in m[#7]
  HD[5299] = 32'b10000101100011000000000000000000;//Loadr m[r[12]] to r[12]
  HD[5300] = 32'b01100001000000000000000000000100;//Load m[#4] to r[8]
  HD[5301] = 32'b10001001100010000000000000000000;//rStore r[12] in m[r[8]]
  HD[5302] = 32'b01100001110000000000000000000111;//Load m[#7] to r[14]
  HD[5303] = 32'b01100001100000000000000000000110;//Load m[#6] to r[12]
  HD[5304] = 32'b10001001110011000000000000000000;//rStore r[14] in m[r[12]]
  HD[5305] = 32'b01100001000000000000000000000100;//Load m[#4] to r[8]
  HD[5306] = 32'b00000101000010000000000000000001;//ADDi r[8], #1 to r[8]
  HD[5307] = 32'b01100101000000000000000000000100;//Store r[8] in m[#4]
  HD[5308] = 32'b01010100000000000000000000010001;//Jump to #17
  HD[5309] = 32'b01100000001000000000000000000000;//Load m[#0] to r[1]
  HD[5310] = 32'b01100000010000000000000000000001;//Load m[#1] to r[2]
  HD[5311] = 32'b01100000011000000000000000000010;//Load m[#2] to r[3]
  HD[5312] = 32'b01100000100000000000000000000011;//Load m[#3] to r[4]
  HD[5313] = 32'b01111000000000000000000000000000;//preio
  HD[5314] = 32'b10000000001000000000000000000000;//Output r[1]
  HD[5315] = 32'b01111000000000000000000000000000;//preio
  HD[5316] = 32'b10000000010000000000000000000000;//Output r[2]
  HD[5317] = 32'b01111000000000000000000000000000;//preio
  HD[5318] = 32'b10000000011000000000000000000000;//Output r[3]
  HD[5319] = 32'b01111000000000000000000000000000;//preio
  HD[5320] = 32'b10000000100000000000000000000000;//Output r[4]
  HD[5321] = 32'b01110000000000000000000000000000;//Hlt
  HD[5322] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]



  //program 7 [line 5440] - Top Down [18]
  HD[5440] = 32'b01101100000000000000000000000000;//Nop
  HD[5441] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[5442] = 32'b01101000001000000100011010100000;//Loadi #18080 to r[1]
  HD[5443] = 32'b01100100001000000000000000000001;//Store r[1] in m[#1]
  HD[5444] = 32'b01101000001000000000000000110010;//Loadi #50 to r[1]
  HD[5445] = 32'b01100100001000000000000000000010;//Store r[1] in m[#2]
  HD[5446] = 32'b01101000001000000000000000000000;//Loadi #0 to r[1]
  HD[5447] = 32'b01100100001000000000000000000100;//Store r[1] in m[#4]
  HD[5448] = 32'b01100000001000000000000000000100;//Load m[#4] to r[1]
  HD[5449] = 32'b01100000010000000000000000000001;//Load m[#1] to r[2]
  HD[5450] = 32'b01011100011000010001000000000000;//SLT if r[1] < r[2], r[3] = 1 else r[3] = 0
  HD[5451] = 32'b01111100000000110000000000000000;//Pre Branch r[3]
  HD[5452] = 32'b01001100000000000000000000001101;//Branch on Zero #13
  HD[5453] = 32'b01101000011000000000000000000010;//Loadi #2 to r[3]
  HD[5454] = 32'b00010100011000100001100000000000;//DIVIDE r[2],r[3] to r[3]
  HD[5455] = 32'b01011100100000010001100000000000;//SLT if r[1] < r[3], r[4] = 1 else r[4] = 0
  HD[5456] = 32'b01011100011000110000100000000000;//SLT if r[3] < r[1], r[3] = 1 else r[3] = 0
  HD[5457] = 32'b00100100011000110010000000000000;//OR r[3],r[4] to r[3]
  HD[5458] = 32'b00110100011000110000000000000000;//NOT r[3] to r[3]
  HD[5459] = 32'b01111100000000110000000000000000;//Pre Branch r[3]
  HD[5460] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[5461] = 32'b01111000000000000000000000000000;//preio
  HD[5462] = 32'b10000000001000000000000000000000;//Output r[1]
  HD[5463] = 32'b01101100000000000000000000000000;//Nop
  HD[5464] = 32'b00000100001000010000000000000001;//ADDi r[1], #1 to r[1]
  HD[5465] = 32'b01010100000000000000000000000111;//Jump to #7
  HD[5466] = 32'b01111000000000000000000000000000;//preio
  HD[5467] = 32'b10000000001000000000000000000000;//Output r[1]
  HD[5468] = 32'b01100000010000000000000000000010;//Load m[#2] to r[2]
  HD[5469] = 32'b01100000001000000000000000000100;//Load m[#4] to r[1]
  HD[5470] = 32'b01011100011000100000100000000000;//SLT if r[2] < r[1], r[3] = 1 else r[3] = 0
  HD[5471] = 32'b01111100000000110000000000000000;//Pre Branch r[3]
  HD[5472] = 32'b01001100000000000000000000001101;//Branch on Zero #13
  HD[5473] = 32'b01101000011000000000000000000010;//Loadi #2 to r[3]
  HD[5474] = 32'b00010000011000100001100000000000;//TIMES r[2],r[3] to r[3]
  HD[5475] = 32'b01011100100000010001100000000000;//SLT if r[1] < r[3], r[4] = 1 else r[4] = 0
  HD[5476] = 32'b01011100011000110000100000000000;//SLT if r[3] < r[1], r[3] = 1 else r[3] = 0
  HD[5477] = 32'b00100100011000110010000000000000;//OR r[3],r[4] to r[3]
  HD[5478] = 32'b00110100011000110000000000000000;//NOT r[3] to r[3]
  HD[5479] = 32'b01111100000000110000000000000000;//Pre Branch r[3]
  HD[5480] = 32'b01001100000000000000000000000011;//Branch on Zero #3
  HD[5481] = 32'b01111000000000000000000000000000;//preio
  HD[5482] = 32'b10000000001000000000000000000000;//Output r[1]
  HD[5483] = 32'b01101100000000000000000000000000;//Nop
  HD[5484] = 32'b00001100001000010000000000000001;//SUBi r[1], #1 to r[1]
  HD[5485] = 32'b01010100000000000000000000011110;//Jump to #30
  HD[5486] = 32'b01111000000000000000000000000000;//preio
  HD[5487] = 32'b10000000001000000000000000000000;//Output r[1]
  HD[5488] = 32'b01110000000000000000000000000000;//Hlt
  HD[5489] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]


  //program 8 [line 5632] - Circle Area [19]
  HD[5632] = 32'b01101100000000000000000000000000;//Nop
  HD[5633] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[5634] = 32'b01101000011000000000110001000110;//Loadi #3142 to r[3]
  HD[5635] = 32'b01111000000000000000000000000000;//preio
  HD[5636] = 32'b01110100101000000000000000000000;//Input to r[5]
  HD[5637] = 32'b00010000101001010010100000000000;//TIMES r[5],r[5] to r[5]
  HD[5638] = 32'b00010000101001010001100000000000;//TIMES r[5],r[3] to r[5]
  HD[5639] = 32'b01101001010000000000001111101000;//Loadi #1000 to r[10]
  HD[5640] = 32'b00010100101001010101000000000000;//DIVIDE r[5],r[10] to r[5]
  HD[5641] = 32'b01111000000000000000000000000000;//preio
  HD[5642] = 32'b10000000101000000000000000000000;//Output r[5]
  HD[5643] = 32'b01110000000000000000000000000000;//Hlt
  HD[5644] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]

  //program 9 [line 5824] - Multiplication [20]
  HD[5824] = 32'b01101100000000000000000000000000;//Nop
  HD[5825] = 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
  HD[5826] = 32'b01111000000000000000000000000000;//preio
  HD[5827] = 32'b01110100001000000000000000000000;//Input to r[1]
  HD[5828] = 32'b01100100001000000000000000000010;//Store r[1] in m[#2]
  HD[5829] = 32'b01111000000000000000000000000000;//preio
  HD[5830] = 32'b01110100001000000000000000000000;//Input to r[1]
  HD[5831] = 32'b01100100001000000000000000000011;//Store r[1] in m[#3]
  HD[5832] = 32'b01100100000000000000000000000100;//Store r[0] in m[#4]
  HD[5833] = 32'b01100000001000000000000000000011;//Load m[#3] to r[1]
  HD[5834] = 32'b01011100100000000000100000000000;//SLT if r[0] < r[1], r[4] = 1 else r[4] = 0
  HD[5835] = 32'b01111100000001000000000000000000;//Pre Branch r[4]
  HD[5836] = 32'b01001100000000000000000000000110;//Branch on Zero #6
  HD[5837] = 32'b01100000110000000000000000000100;//Load m[#4] to r[6]
  HD[5838] = 32'b01100000111000000000000000000010;//Load m[#2] to r[7]
  HD[5839] = 32'b00000000111001100011100000000000;//ADD r[6],r[7] to r[7]
  HD[5840] = 32'b01100100111000000000000000000100;//Store r[7] in m[#4]
  HD[5841] = 32'b00001100001000010000000000000001;//SUBi r[1], #1 to r[1]
  HD[5842] = 32'b01010100000000000000000000001010;//Jump to #10
  HD[5843] = 32'b01100001010000000000000000000100;//Load m[#4] to r[10]
  HD[5844] = 32'b01111000000000000000000000000000;//preio
  HD[5845] = 32'b10000001010000000000000000000000;//Output r[10]
  HD[5846] = 32'b01110000000000000000000000000000;//Hlt
  HD[5847] = 32'b00000000000000000000000000000000;//ADD r[0],r[0] to r[0]


end


    always @ (posedge clock)
    begin
      // Write
      if (flag_write_hd)
        HD[hd_address] <= data_write;

      hd_local_address <= hd_address;
    //  sector_address <= sector;
    end


	// Continuous assignment implies read returns NEW data.
	// This is the natural behavior of the TriMatrix memory
	// blocks in Single Port mode.
	assign output_hard_drive = HD[hd_local_address];

endmodule
